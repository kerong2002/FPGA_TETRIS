
module IMG(
    input wire [9:0] x,
    input wire [9:0] y,
    output reg [23:0] pixel
);

        always @(*) begin
        case (y)
            10'd0: case (x)
                10'd0: pixel <= 24'h22_41_81;
                10'd1: pixel <= 24'h43_87_FF;
                10'd2: pixel <= 24'h85_FF_1F;
                10'd3: pixel <= 24'hFF_20_43;
                10'd4: pixel <= 24'h20_43_87;
                10'd5: pixel <= 24'h1C_49_FF;
                10'd6: pixel <= 24'h38_FF_08;
                10'd7: pixel <= 24'hFF_0B_18;
                10'd8: pixel <= 24'h0B_18_38;
                10'd9: pixel <= 24'h18_38_FF;
                10'd10: pixel <= 24'h38_FF_0B;
                10'd11: pixel <= 24'hFF_0B_18;
                10'd12: pixel <= 24'h0B_18_38;
                10'd13: pixel <= 24'h18_38_FF;
                10'd14: pixel <= 24'h33_FF_0B;
                10'd15: pixel <= 24'hFF_0F_12;
                10'd16: pixel <= 24'hEB_25_3D;
                10'd17: pixel <= 24'h4A_65_FF;
                10'd18: pixel <= 24'h67_FF_F0;
                10'd19: pixel <= 24'hFF_EF_4B;
                10'd20: pixel <= 24'hEF_4B_67;
                10'd21: pixel <= 24'h4B_67_FF;
                10'd22: pixel <= 24'h38_FF_EF;
                10'd23: pixel <= 24'hFF_EE_2A;
                10'd24: pixel <= 24'h0B_18_38;
                10'd25: pixel <= 24'h17_38_FF;
                10'd26: pixel <= 24'h38_FF_0C;
                10'd27: pixel <= 24'hFF_0C_17;
                10'd28: pixel <= 24'h0B_18_38;
                10'd29: pixel <= 24'h16_38_FF;
                10'd30: pixel <= 24'h1E_FF_09;
                10'd31: pixel <= 24'hFF_EF_88;
                10'd32: pixel <= 24'hFC_CA_21;
                10'd33: pixel <= 24'hCA_21_FF;
                10'd34: pixel <= 24'h21_FF_FE;
                10'd35: pixel <= 24'hFF_FE_CA;
                10'd36: pixel <= 24'hFF_CB_22;
                10'd37: pixel <= 24'hCB_22_FF;
                10'd38: pixel <= 24'h22_FF_FF;
                10'd39: pixel <= 24'hFF_FF_CB;
                10'd40: pixel <= 24'hFF_CB_22;
                10'd41: pixel <= 24'hCB_22_FF;
                10'd42: pixel <= 24'h22_FF_FF;
                10'd43: pixel <= 24'hFF_FF_CB;
                10'd44: pixel <= 24'hFB_CA_25;
                10'd45: pixel <= 24'h69_25_FF;
                10'd46: pixel <= 24'h38_FF_F2;
                10'd47: pixel <= 24'hFF_0B_18;
                10'd48: pixel <= 24'h0C_19_39;
                10'd49: pixel <= 24'h18_38_FF;
                10'd50: pixel <= 24'h38_FF_0B;
                10'd51: pixel <= 24'hFF_0B_18;
                10'd52: pixel <= 24'h0B_18_38;
                10'd53: pixel <= 24'h18_38_FF;
                10'd54: pixel <= 24'h38_FF_0B;
                10'd55: pixel <= 24'hFF_0B_18;
                10'd56: pixel <= 24'h0A_0C_0E;
                10'd57: pixel <= 24'hBA_15_FF;
                10'd58: pixel <= 24'h21_FF_F3;
                10'd59: pixel <= 24'hFF_FB_E1;
                10'd60: pixel <= 24'hFB_E1_21;
                10'd61: pixel <= 24'hE1_21_FF;
                10'd62: pixel <= 24'h1F_FF_FB;
                10'd63: pixel <= 24'hFF_FB_E1;
                10'd64: pixel <= 24'hE8_AA_3D;
                10'd65: pixel <= 24'h18_38_FF;
                10'd66: pixel <= 24'h38_FF_09;
                10'd67: pixel <= 24'hFF_0B_18;
                10'd68: pixel <= 24'h0B_18_38;
                10'd69: pixel <= 24'h18_38_FF;
                10'd70: pixel <= 24'h38_FF_0B;
                10'd71: pixel <= 24'hFF_0B_18;
                10'd72: pixel <= 24'h55_B0_44;
                10'd73: pixel <= 24'hC5_4D_FF;
                10'd74: pixel <= 24'h4C_FF_90;
                10'd75: pixel <= 24'hFF_8F_C8;
                10'd76: pixel <= 24'h8F_C8_4C;
                10'd77: pixel <= 24'hC8_4C_FF;
                10'd78: pixel <= 24'h49_FF_8F;
                10'd79: pixel <= 24'hFF_49_B1;
                10'd80: pixel <= 24'h43_B2_46;
                10'd81: pixel <= 24'hC8_4C_FF;
                10'd82: pixel <= 24'h4C_FF_91;
                10'd83: pixel <= 24'hFF_91_C7;
                10'd84: pixel <= 24'h8F_C8_4C;
                10'd85: pixel <= 24'hC8_4C_FF;
                10'd86: pixel <= 24'h4D_FF_8F;
                10'd87: pixel <= 24'hFF_90_C9;
                10'd88: pixel <= 24'h3C_B0_4B;
                10'd89: pixel <= 24'h1A_33_FF;
                10'd90: pixel <= 24'h34_FF_06;
                10'd91: pixel <= 24'hFF_09_17;
                10'd92: pixel <= 24'h0B_18_38;
                10'd93: pixel <= 24'h18_38_FF;
                10'd94: pixel <= 24'hD3_FF_0B;
                10'd95: pixel <= 24'hFF_07_A0;
                10'd96: pixel <= 24'h6B_CD_DB;
                10'd97: pixel <= 24'hCC_DB_FF;
                10'd98: pixel <= 24'hDB_FF_6C;
                10'd99: pixel <= 24'hFF_6C_CC;
            endcase
            10'd1: case (x)
                10'd0: pixel <= 24'hFD_D0_22;
                10'd1: pixel <= 24'hD0_24_FF;
                10'd2: pixel <= 24'h22_FF_FD;
                10'd3: pixel <= 24'hFF_FD_D0;
                10'd4: pixel <= 24'hFD_D0_22;
                10'd5: pixel <= 24'hD0_22_FF;
                10'd6: pixel <= 24'h22_FF_FD;
                10'd7: pixel <= 24'hFF_FD_D0;
                10'd8: pixel <= 24'hFB_CE_23;
                10'd9: pixel <= 24'hD0_1F_FF;
                10'd10: pixel <= 24'h1E_FF_FA;
                10'd11: pixel <= 24'hFF_E9_70;
                10'd12: pixel <= 24'h18_0A_17;
                10'd13: pixel <= 24'h18_38_FF;
                10'd14: pixel <= 24'h3A_FF_09;
                10'd15: pixel <= 24'hFF_0B_17;
                10'd16: pixel <= 24'h0B_17_3A;
                10'd17: pixel <= 24'h17_3A_FF;
                10'd18: pixel <= 24'h3A_FF_0B;
                10'd19: pixel <= 24'hFF_0B_17;
                10'd20: pixel <= 24'h0B_17_3A;
                10'd21: pixel <= 24'h17_3A_FF;
                10'd22: pixel <= 24'h12_FF_0B;
                10'd23: pixel <= 24'hFF_0A_0B;
                10'd24: pixel <= 24'hFE_B6_23;
                10'd25: pixel <= 24'h87_1D_FF;
                10'd26: pixel <= 24'h1C_FF_F3;
                10'd27: pixel <= 24'hFF_F4_88;
                10'd28: pixel <= 24'hF2_81_1C;
                10'd29: pixel <= 24'h86_1B_FF;
                10'd30: pixel <= 24'h3E_FF_F1;
                10'd31: pixel <= 24'hFF_E7_A8;
                10'd32: pixel <= 24'h09_18_3A;
                10'd33: pixel <= 24'h17_3A_FF;
                10'd34: pixel <= 24'h3A_FF_0B;
                10'd35: pixel <= 24'hFF_0B_17;
                10'd36: pixel <= 24'h0B_17_3A;
                10'd37: pixel <= 24'h17_3A_FF;
                10'd38: pixel <= 24'h44_FF_0B;
                10'd39: pixel <= 24'hFF_54_AE;
                10'd40: pixel <= 24'h17_71_38;
                10'd41: pixel <= 24'h72_2F_FF;
                10'd42: pixel <= 24'h30_FF_18;
                10'd43: pixel <= 24'hFF_1C_73;
                10'd44: pixel <= 24'h27_7C_2B;
                10'd45: pixel <= 24'hB2_46_FF;
                10'd46: pixel <= 24'h49_FF_48;
                10'd47: pixel <= 24'hFF_46_B3;
                10'd48: pixel <= 24'h88_CE_64;
                10'd49: pixel <= 24'hCB_4C_FF;
                10'd50: pixel <= 24'h4E_FF_90;
                10'd51: pixel <= 24'hFF_93_C9;
                10'd52: pixel <= 24'h93_C9_52;
                10'd53: pixel <= 24'hC9_4E_FF;
                10'd54: pixel <= 24'h44_FF_95;
                10'd55: pixel <= 24'hFF_31_A3;
                10'd56: pixel <= 24'h0C_16_3A;
                10'd57: pixel <= 24'h17_38_FF;
                10'd58: pixel <= 24'h3A_FF_0C;
                10'd59: pixel <= 24'hFF_0B_17;
                10'd60: pixel <= 24'h0B_17_3A;
                10'd61: pixel <= 24'hA1_D4_FF;
                10'd62: pixel <= 24'hDB_FF_08;
                10'd63: pixel <= 24'hFF_6C_CC;
                10'd64: pixel <= 24'h6F_CE_DE;
                10'd65: pixel <= 24'hCD_DD_FF;
                10'd66: pixel <= 24'hDD_FF_6E;
                10'd67: pixel <= 24'hFF_70_CA;
                10'd68: pixel <= 24'h11_7D_BF;
                10'd69: pixel <= 24'h17_38_FF;
                10'd70: pixel <= 24'h3A_FF_0C;
                10'd71: pixel <= 24'hFF_0B_17;
                10'd72: pixel <= 24'h0B_17_3A;
                10'd73: pixel <= 24'h13_3E_FF;
                10'd74: pixel <= 24'h8A_FF_12;
                10'd75: pixel <= 24'hFF_9C_2B;
                10'd76: pixel <= 24'hBC_59_A3;
                10'd77: pixel <= 24'h59_A1_FF;
                10'd78: pixel <= 24'hA1_FF_BC;
                10'd79: pixel <= 24'hFF_BC_59;
                10'd80: pixel <= 24'hBC_59_A1;
                10'd81: pixel <= 24'h58_A0_FF;
                10'd82: pixel <= 24'h8B_FF_BA;
                10'd83: pixel <= 24'hFF_92_28;
                10'd84: pixel <= 24'h12_1A_3F;
                10'd85: pixel <= 24'h17_3C_FF;
                10'd86: pixel <= 24'h3A_FF_0B;
                10'd87: pixel <= 24'hFF_0B_17;
                10'd88: pixel <= 24'h0B_17_3A;
                10'd89: pixel <= 24'h17_3A_FF;
                10'd90: pixel <= 24'h3A_FF_0B;
                10'd91: pixel <= 24'hFF_0B_17;
                10'd92: pixel <= 24'h0B_17_3A;
                10'd93: pixel <= 24'h17_3A_FF;
                10'd94: pixel <= 24'h85_FF_0B;
                10'd95: pixel <= 24'hFF_20_43;
                10'd96: pixel <= 24'h20_45_88;
                10'd97: pixel <= 24'h44_8A_FF;
                10'd98: pixel <= 24'h81_FF_20;
                10'd99: pixel <= 24'hFF_21_41;
            endcase
            10'd2: case (x)
                10'd0: pixel <= 24'h0C_18_3D;
                10'd1: pixel <= 24'h18_3D_FF;
                10'd2: pixel <= 24'h3D_FF_0C;
                10'd3: pixel <= 24'hFF_0C_18;
                10'd4: pixel <= 24'h0C_18_3D;
                10'd5: pixel <= 24'hB0_42_FF;
                10'd6: pixel <= 24'h3B_FF_51;
                10'd7: pixel <= 24'hFF_15_75;
                10'd8: pixel <= 24'h12_76_3D;
                10'd9: pixel <= 24'h76_3B_FF;
                10'd10: pixel <= 24'h3D_FF_13;
                10'd11: pixel <= 24'hFF_15_74;
                10'd12: pixel <= 24'h48_B1_4B;
                10'd13: pixel <= 24'h40_3C_FF;
                10'd14: pixel <= 24'h47_FF_1D;
                10'd15: pixel <= 24'hFF_39_B0;
                10'd16: pixel <= 24'h14_75_45;
                10'd17: pixel <= 24'h76_3B_FF;
                10'd18: pixel <= 24'h3B_FF_13;
                10'd19: pixel <= 24'hFF_13_76;
                10'd20: pixel <= 24'h14_77_3C;
                10'd21: pixel <= 24'h8C_40_FF;
                10'd22: pixel <= 24'h50_FF_24;
                10'd23: pixel <= 24'hFF_31_85;
                10'd24: pixel <= 24'h0C_17_38;
                10'd25: pixel <= 24'h18_3D_FF;
                10'd26: pixel <= 24'h3C_FF_0C;
                10'd27: pixel <= 24'hFF_0B_17;
                10'd28: pixel <= 24'h08_A2_D2;
                10'd29: pixel <= 24'hCB_DD_FF;
                10'd30: pixel <= 24'hDB_FF_6E;
                10'd31: pixel <= 24'hFF_6B_CD;
                10'd32: pixel <= 24'h6E_CB_DB;
                10'd33: pixel <= 24'hC9_DC_FF;
                10'd34: pixel <= 24'hBF_FF_6E;
                10'd35: pixel <= 24'hFF_11_7D;
                10'd36: pixel <= 24'h0D_18_39;
                10'd37: pixel <= 24'h18_3D_FF;
                10'd38: pixel <= 24'h3D_FF_0C;
                10'd39: pixel <= 24'hFF_0C_18;
                10'd40: pixel <= 24'h0C_18_3B;
                10'd41: pixel <= 24'h39_7B_FF;
                10'd42: pixel <= 24'h8D_FF_6E;
                10'd43: pixel <= 24'hFF_A0_2C;
                10'd44: pixel <= 24'hBC_59_A1;
                10'd45: pixel <= 24'h59_A1_FF;
                10'd46: pixel <= 24'hA2_FF_BC;
                10'd47: pixel <= 24'hFF_BD_5B;
                10'd48: pixel <= 24'hBD_5B_A2;
                10'd49: pixel <= 24'h58_AB_FF;
                10'd50: pixel <= 24'h78_FF_BD;
                10'd51: pixel <= 24'hFF_7C_2A;
                10'd52: pixel <= 24'h0B_16_3E;
                10'd53: pixel <= 24'h17_3C_FF;
                10'd54: pixel <= 24'h3D_FF_0B;
                10'd55: pixel <= 24'hFF_0C_18;
                10'd56: pixel <= 24'h0C_18_3D;
                10'd57: pixel <= 24'h18_3D_FF;
                10'd58: pixel <= 24'h3D_FF_0C;
                10'd59: pixel <= 24'hFF_0C_18;
                10'd60: pixel <= 24'h0C_18_3B;
                10'd61: pixel <= 24'h45_89_FF;
                10'd62: pixel <= 24'h8A_FF_22;
                10'd63: pixel <= 24'hFF_22_47;
                10'd64: pixel <= 24'h25_45_8A;
                10'd65: pixel <= 24'h40_83_FF;
                10'd66: pixel <= 24'h81_FF_22;
                10'd67: pixel <= 24'hFF_22_41;
                10'd68: pixel <= 24'h20_45_88;
                10'd69: pixel <= 24'h45_88_FF;
                10'd70: pixel <= 24'h88_FF_20;
                10'd71: pixel <= 24'hFF_23_43;
                10'd72: pixel <= 24'h09_1D_4A;
                10'd73: pixel <= 24'h17_3A_FF;
                10'd74: pixel <= 24'h3A_FF_0B;
                10'd75: pixel <= 24'hFF_0B_17;
                10'd76: pixel <= 24'h0B_17_3A;
                10'd77: pixel <= 24'h17_3A_FF;
                10'd78: pixel <= 24'h3A_FF_0B;
                10'd79: pixel <= 24'hFF_0B_17;
                10'd80: pixel <= 24'h0B_17_3A;
                10'd81: pixel <= 24'h12_35_FF;
                10'd82: pixel <= 24'h41_FF_0F;
                10'd83: pixel <= 24'hFF_EB_25;
                10'd84: pixel <= 24'hF0_4A_67;
                10'd85: pixel <= 24'h4B_67_FF;
                10'd86: pixel <= 24'h67_FF_EF;
                10'd87: pixel <= 24'hFF_EF_4B;
                10'd88: pixel <= 24'hEF_4B_67;
                10'd89: pixel <= 24'h2A_38_FF;
                10'd90: pixel <= 24'h3A_FF_EE;
                10'd91: pixel <= 24'hFF_0B_17;
                10'd92: pixel <= 24'h0B_17_3A;
                10'd93: pixel <= 24'h17_3A_FF;
                10'd94: pixel <= 24'h3A_FF_0B;
                10'd95: pixel <= 24'hFF_0B_17;
                10'd96: pixel <= 24'h09_16_3A;
                10'd97: pixel <= 24'h87_1F_FF;
                10'd98: pixel <= 24'h21_FF_EE;
                10'd99: pixel <= 24'hFF_FD_CE;
            endcase
            10'd3: case (x)
                10'd0: pixel <= 24'h74_CF_E9;
                10'd1: pixel <= 24'h7F_BA_FF;
                10'd2: pixel <= 24'h3E_FF_12;
                10'd3: pixel <= 24'hFF_0E_18;
                10'd4: pixel <= 24'h0D_19_3E;
                10'd5: pixel <= 24'h18_3E_FF;
                10'd6: pixel <= 24'h3E_FF_0E;
                10'd7: pixel <= 24'hFF_0E_18;
                10'd8: pixel <= 24'h0D_19_3C;
                10'd9: pixel <= 24'h3F_96_FF;
                10'd10: pixel <= 24'hA8_FF_A3;
                10'd11: pixel <= 24'hFF_C0_58;
                10'd12: pixel <= 24'hBB_5C_A0;
                10'd13: pixel <= 24'h5B_A2_FF;
                10'd14: pixel <= 24'hA2_FF_BD;
                10'd15: pixel <= 24'hFF_BD_5B;
                10'd16: pixel <= 24'hBD_5B_A0;
                10'd17: pixel <= 24'h31_8A_FF;
                10'd18: pixel <= 24'h67_FF_9C;
                10'd19: pixel <= 24'hFF_66_26;
                10'd20: pixel <= 24'h0D_17_3D;
                10'd21: pixel <= 24'h19_3E_FF;
                10'd22: pixel <= 24'h3E_FF_0D;
                10'd23: pixel <= 24'hFF_0D_19;
                10'd24: pixel <= 24'h0E_18_3E;
                10'd25: pixel <= 24'h19_3E_FF;
                10'd26: pixel <= 24'h3D_FF_0D;
                10'd27: pixel <= 24'hFF_0C_18;
                10'd28: pixel <= 24'h24_46_8A;
                10'd29: pixel <= 24'h48_8D_FF;
                10'd30: pixel <= 24'h8C_FF_23;
                10'd31: pixel <= 24'hFF_23_4A;
                10'd32: pixel <= 24'h22_41_81;
                10'd33: pixel <= 24'h3F_83_FF;
                10'd34: pixel <= 24'h8A_FF_24;
                10'd35: pixel <= 24'hFF_22_47;
                10'd36: pixel <= 24'h22_47_8A;
                10'd37: pixel <= 24'h47_8A_FF;
                10'd38: pixel <= 24'h49_FF_22;
                10'd39: pixel <= 24'hFF_08_1C;
                10'd40: pixel <= 24'h0C_18_3B;
                10'd41: pixel <= 24'h18_3D_FF;
                10'd42: pixel <= 24'h3D_FF_0C;
                10'd43: pixel <= 24'hFF_0C_18;
                10'd44: pixel <= 24'h0C_18_3D;
                10'd45: pixel <= 24'h18_3D_FF;
                10'd46: pixel <= 24'h3D_FF_0C;
                10'd47: pixel <= 24'hFF_0C_18;
                10'd48: pixel <= 24'h0D_12_37;
                10'd49: pixel <= 24'h26_3F_FF;
                10'd50: pixel <= 24'h65_FF_E9;
                10'd51: pixel <= 24'hFF_F0_4A;
                10'd52: pixel <= 24'hEF_4B_67;
                10'd53: pixel <= 24'h4B_67_FF;
                10'd54: pixel <= 24'h67_FF_EF;
                10'd55: pixel <= 24'hFF_EF_4B;
                10'd56: pixel <= 24'hEE_2A_3A;
                10'd57: pixel <= 24'h18_3D_FF;
                10'd58: pixel <= 24'h3D_FF_0C;
                10'd59: pixel <= 24'hFF_0C_18;
                10'd60: pixel <= 24'h0C_18_3D;
                10'd61: pixel <= 24'h18_3D_FF;
                10'd62: pixel <= 24'h3C_FF_0C;
                10'd63: pixel <= 24'hFF_0B_17;
                10'd64: pixel <= 24'hF1_87_20;
                10'd65: pixel <= 24'hD3_23_FF;
                10'd66: pixel <= 24'h24_FF_FA;
                10'd67: pixel <= 24'hFF_FD_D3;
                10'd68: pixel <= 24'hFA_D5_22;
                10'd69: pixel <= 24'hD3_22_FF;
                10'd70: pixel <= 24'h20_FF_FD;
                10'd71: pixel <= 24'hFF_F6_D4;
                10'd72: pixel <= 24'hFF_D1_2F;
                10'd73: pixel <= 24'hBC_35_FF;
                10'd74: pixel <= 24'h14_FF_FF;
                10'd75: pixel <= 24'hFF_DE_5D;
                10'd76: pixel <= 24'hDA_2C_13;
                10'd77: pixel <= 24'h6E_25_FF;
                10'd78: pixel <= 24'h3C_FF_EB;
                10'd79: pixel <= 24'hFF_0B_17;
                10'd80: pixel <= 24'h09_18_3C;
                10'd81: pixel <= 24'h17_3C_FF;
                10'd82: pixel <= 24'h3B_FF_0B;
                10'd83: pixel <= 24'hFF_0C_18;
                10'd84: pixel <= 24'h0C_18_3D;
                10'd85: pixel <= 24'h18_3D_FF;
                10'd86: pixel <= 24'h3D_FF_0C;
                10'd87: pixel <= 24'hFF_0C_18;
                10'd88: pixel <= 24'h0C_18_3D;
                10'd89: pixel <= 24'h0E_11_FF;
                10'd90: pixel <= 24'h21_FF_0A;
                10'd91: pixel <= 24'hFF_FF_B4;
                10'd92: pixel <= 24'hF9_86_1D;
                10'd93: pixel <= 24'h87_1F_FF;
                10'd94: pixel <= 24'h1F_FF_F5;
                10'd95: pixel <= 24'hFF_F5_87;
                10'd96: pixel <= 24'hF4_86_1E;
                10'd97: pixel <= 24'hAA_41_FF;
                10'd98: pixel <= 24'h3D_FF_E6;
                10'd99: pixel <= 24'hFF_0C_18;
            endcase
            10'd4: case (x)
                10'd0: pixel <= 24'h24_3F_83;
                10'd1: pixel <= 24'h49_8E_FF;
                10'd2: pixel <= 24'h8C_FF_24;
                10'd3: pixel <= 24'hFF_23_4A;
                10'd4: pixel <= 24'h22_47_8A;
                10'd5: pixel <= 24'h1E_4C_FF;
                10'd6: pixel <= 24'h3E_FF_0A;
                10'd7: pixel <= 24'hFF_0D_19;
                10'd8: pixel <= 24'h0D_19_3E;
                10'd9: pixel <= 24'h19_3E_FF;
                10'd10: pixel <= 24'h3E_FF_0D;
                10'd11: pixel <= 24'hFF_0E_18;
                10'd12: pixel <= 24'h0D_19_3E;
                10'd13: pixel <= 24'h18_3E_FF;
                10'd14: pixel <= 24'h3B_FF_0E;
                10'd15: pixel <= 24'hFF_12_15;
                10'd16: pixel <= 24'hEB_25_3D;
                10'd17: pixel <= 24'h4A_65_FF;
                10'd18: pixel <= 24'h67_FF_F0;
                10'd19: pixel <= 24'hFF_EF_4B;
                10'd20: pixel <= 24'hEF_4B_67;
                10'd21: pixel <= 24'h4B_67_FF;
                10'd22: pixel <= 24'h38_FF_EF;
                10'd23: pixel <= 24'hFF_EE_2A;
                10'd24: pixel <= 24'h0E_18_3E;
                10'd25: pixel <= 24'h19_3E_FF;
                10'd26: pixel <= 24'h3E_FF_0D;
                10'd27: pixel <= 24'hFF_0D_19;
                10'd28: pixel <= 24'h0D_19_3E;
                10'd29: pixel <= 24'h17_41_FF;
                10'd30: pixel <= 24'h1A_FF_0C;
                10'd31: pixel <= 24'hFF_EF_83;
                10'd32: pixel <= 24'hFF_D4_40;
                10'd33: pixel <= 24'h5F_1D_FF;
                10'd34: pixel <= 24'h1C_FF_EB;
                10'd35: pixel <= 24'hFF_E2_32;
                10'd36: pixel <= 24'hED_2B_24;
                10'd37: pixel <= 24'h29_26_FF;
                10'd38: pixel <= 24'h26_FF_EC;
                10'd39: pixel <= 24'hFF_ED_2A;
                10'd40: pixel <= 24'hEB_2A_24;
                10'd41: pixel <= 24'h2C_24_FF;
                10'd42: pixel <= 24'h25_FF_EC;
                10'd43: pixel <= 24'hFF_F5_6C;
                10'd44: pixel <= 24'h14_17_37;
                10'd45: pixel <= 24'h19_3E_FF;
                10'd46: pixel <= 24'h40_FF_0D;
                10'd47: pixel <= 24'hFF_0E_18;
                10'd48: pixel <= 24'h0E_18_40;
                10'd49: pixel <= 24'h19_3E_FF;
                10'd50: pixel <= 24'h3E_FF_0D;
                10'd51: pixel <= 24'hFF_0D_19;
                10'd52: pixel <= 24'h0E_18_3E;
                10'd53: pixel <= 24'h19_3E_FF;
                10'd54: pixel <= 24'h3E_FF_0D;
                10'd55: pixel <= 24'hFF_0D_19;
                10'd56: pixel <= 24'h0B_0F_12;
                10'd57: pixel <= 24'hB3_20_FF;
                10'd58: pixel <= 24'h20_FF_FF;
                10'd59: pixel <= 24'hFF_F5_89;
                10'd60: pixel <= 24'hF7_88_20;
                10'd61: pixel <= 24'h89_1E_FF;
                10'd62: pixel <= 24'h1F_FF_F5;
                10'd63: pixel <= 24'hFF_F5_87;
                10'd64: pixel <= 24'hE6_AA_41;
                10'd65: pixel <= 24'h18_3E_FF;
                10'd66: pixel <= 24'h3E_FF_0E;
                10'd67: pixel <= 24'hFF_0D_19;
                10'd68: pixel <= 24'h0D_19_3E;
                10'd69: pixel <= 24'h19_3E_FF;
                10'd70: pixel <= 24'h3E_FF_0D;
                10'd71: pixel <= 24'hFF_0D_19;
                10'd72: pixel <= 24'h52_AF_42;
                10'd73: pixel <= 24'h79_3F_FF;
                10'd74: pixel <= 24'h3E_FF_17;
                10'd75: pixel <= 24'hFF_14_79;
                10'd76: pixel <= 24'h14_79_3E;
                10'd77: pixel <= 24'h78_3E_FF;
                10'd78: pixel <= 24'h4B_FF_16;
                10'd79: pixel <= 24'hFF_48_B1;
                10'd80: pixel <= 24'h0E_19_3C;
                10'd81: pixel <= 24'hB0_4B_FF;
                10'd82: pixel <= 24'h34_FF_42;
                10'd83: pixel <= 24'hFF_11_76;
                10'd84: pixel <= 24'h16_78_3C;
                10'd85: pixel <= 24'h7A_3F_FF;
                10'd86: pixel <= 24'h3F_FF_15;
                10'd87: pixel <= 24'hFF_15_7A;
                10'd88: pixel <= 24'h14_79_3A;
                10'd89: pixel <= 24'hAE_53_FF;
                10'd90: pixel <= 24'h38_FF_43;
                10'd91: pixel <= 24'hFF_0A_1B;
                10'd92: pixel <= 24'h0B_1A_3C;
                10'd93: pixel <= 24'h19_3E_FF;
                10'd94: pixel <= 24'hD5_FF_0D;
                10'd95: pixel <= 24'hFF_07_A0;
                10'd96: pixel <= 24'h26_5E_AD;
                10'd97: pixel <= 24'h60_A6_FF;
                10'd98: pixel <= 24'hB6_FF_22;
                10'd99: pixel <= 24'hFF_38_7B;
            endcase
            10'd5: case (x)
                10'd0: pixel <= 24'hED_2F_26;
                10'd1: pixel <= 24'h2D_23_FF;
                10'd2: pixel <= 24'h27_FF_ED;
                10'd3: pixel <= 24'hFF_EB_2D;
                10'd4: pixel <= 24'hF0_76_1D;
                10'd5: pixel <= 24'h9C_3A_FF;
                10'd6: pixel <= 24'h39_FF_EB;
                10'd7: pixel <= 24'hFF_E9_93;
                10'd8: pixel <= 24'hEC_8B_33;
                10'd9: pixel <= 24'h84_4F_FF;
                10'd10: pixel <= 24'h40_FF_D7;
                10'd11: pixel <= 24'hFF_0E_18;
                10'd12: pixel <= 24'h0E_1A_3F;
                10'd13: pixel <= 24'h19_41_FF;
                10'd14: pixel <= 24'h41_FF_10;
                10'd15: pixel <= 24'hFF_10_19;
                10'd16: pixel <= 24'h0E_1A_3F;
                10'd17: pixel <= 24'h1A_3F_FF;
                10'd18: pixel <= 24'h3F_FF_0E;
                10'd19: pixel <= 24'hFF_10_19;
                10'd20: pixel <= 24'h0E_1A_3F;
                10'd21: pixel <= 24'h1A_3F_FF;
                10'd22: pixel <= 24'h13_FF_0E;
                10'd23: pixel <= 24'hFF_0E_0F;
                10'd24: pixel <= 24'hFF_B3_20;
                10'd25: pixel <= 24'h8A_20_FF;
                10'd26: pixel <= 24'h20_FF_F3;
                10'd27: pixel <= 24'hFF_F7_88;
                10'd28: pixel <= 24'hF5_89_1E;
                10'd29: pixel <= 24'h88_1D_FF;
                10'd30: pixel <= 24'h41_FF_F4;
                10'd31: pixel <= 24'hFF_E8_A9;
                10'd32: pixel <= 24'h10_19_3F;
                10'd33: pixel <= 24'h1A_3F_FF;
                10'd34: pixel <= 24'h3F_FF_0E;
                10'd35: pixel <= 24'hFF_0E_1A;
                10'd36: pixel <= 24'h0E_1A_3F;
                10'd37: pixel <= 24'h1A_3F_FF;
                10'd38: pixel <= 24'h44_FF_0E;
                10'd39: pixel <= 24'hFF_54_B0;
                10'd40: pixel <= 24'h16_7B_40;
                10'd41: pixel <= 24'h7A_3F_FF;
                10'd42: pixel <= 24'h3F_FF_15;
                10'd43: pixel <= 24'hFF_14_7B;
                10'd44: pixel <= 24'h15_7A_3D;
                10'd45: pixel <= 24'hAF_48_FF;
                10'd46: pixel <= 24'h42_FF_48;
                10'd47: pixel <= 24'hFF_11_1A;
                10'd48: pixel <= 24'h0A_1B_39;
                10'd49: pixel <= 24'hB0_53_FF;
                10'd50: pixel <= 24'h40_FF_3F;
                10'd51: pixel <= 24'hFF_16_7B;
                10'd52: pixel <= 24'h14_7B_3F;
                10'd53: pixel <= 24'h7A_3F_FF;
                10'd54: pixel <= 24'h3F_FF_15;
                10'd55: pixel <= 24'hFF_15_7A;
                10'd56: pixel <= 24'h11_7B_3C;
                10'd57: pixel <= 24'h84_3B_FF;
                10'd58: pixel <= 24'h43_FF_1D;
                10'd59: pixel <= 24'hFF_0E_19;
                10'd60: pixel <= 24'h10_19_41;
                10'd61: pixel <= 24'hA2_D6_FF;
                10'd62: pixel <= 24'hAF_FF_06;
                10'd63: pixel <= 24'hFF_27_61;
                10'd64: pixel <= 24'h27_62_AB;
                10'd65: pixel <= 24'h63_AD_FF;
                10'd66: pixel <= 24'hAB_FF_24;
                10'd67: pixel <= 24'hFF_25_62;
                10'd68: pixel <= 24'h13_7F_C1;
                10'd69: pixel <= 24'h19_43_FF;
                10'd70: pixel <= 24'h3F_FF_10;
                10'd71: pixel <= 24'hFF_0E_1A;
                10'd72: pixel <= 24'h10_19_3F;
                10'd73: pixel <= 24'h19_3F_FF;
                10'd74: pixel <= 24'h3F_FF_10;
                10'd75: pixel <= 24'hFF_10_19;
                10'd76: pixel <= 24'h10_1C_43;
                10'd77: pixel <= 24'h32_92_FF;
                10'd78: pixel <= 24'hA5_FF_9A;
                10'd79: pixel <= 24'hFF_C0_60;
                10'd80: pixel <= 24'hBD_5B_A2;
                10'd81: pixel <= 24'h5B_A2_FF;
                10'd82: pixel <= 24'hA2_FF_BD;
                10'd83: pixel <= 24'hFF_BD_5B;
                10'd84: pixel <= 24'hBD_5A_A4;
                10'd85: pixel <= 24'h2E_92_FF;
                10'd86: pixel <= 24'h3D_FF_A1;
                10'd87: pixel <= 24'hFF_18_15;
                10'd88: pixel <= 24'h0E_1A_3F;
                10'd89: pixel <= 24'h1A_3F_FF;
                10'd90: pixel <= 24'h3F_FF_0E;
                10'd91: pixel <= 24'hFF_10_19;
                10'd92: pixel <= 24'h0E_1A_3F;
                10'd93: pixel <= 24'h18_3D_FF;
                10'd94: pixel <= 24'h8B_FF_0C;
                10'd95: pixel <= 24'hFF_25_47;
                10'd96: pixel <= 24'h24_49_8E;
                10'd97: pixel <= 24'h4A_8E_FF;
                10'd98: pixel <= 24'h81_FF_23;
                10'd99: pixel <= 24'hFF_22_41;
            endcase
            10'd6: case (x)
                10'd0: pixel <= 24'h0F_1B_42;
                10'd1: pixel <= 24'h1A_42_FF;
                10'd2: pixel <= 24'h42_FF_11;
                10'd3: pixel <= 24'hFF_11_1A;
                10'd4: pixel <= 24'h11_1A_42;
                10'd5: pixel <= 24'hAF_42_FF;
                10'd6: pixel <= 24'h42_FF_52;
                10'd7: pixel <= 24'hFF_17_7E;
                10'd8: pixel <= 24'h17_7E_42;
                10'd9: pixel <= 24'h7F_40_FF;
                10'd10: pixel <= 24'h3E_FF_17;
                10'd11: pixel <= 24'hFF_19_7E;
                10'd12: pixel <= 24'h49_B1_49;
                10'd13: pixel <= 24'h1B_43_FF;
                10'd14: pixel <= 24'h40_FF_12;
                10'd15: pixel <= 24'hFF_12_1A;
                10'd16: pixel <= 24'h54_AA_66;
                10'd17: pixel <= 24'h9B_47_FF;
                10'd18: pixel <= 24'h40_FF_2E;
                10'd19: pixel <= 24'hFF_17_7F;
                10'd20: pixel <= 24'h17_7D_3F;
                10'd21: pixel <= 24'h7D_3F_FF;
                10'd22: pixel <= 24'h44_FF_16;
                10'd23: pixel <= 24'hFF_15_7F;
                10'd24: pixel <= 24'h42_B4_53;
                10'd25: pixel <= 24'h36_39_FF;
                10'd26: pixel <= 24'h42_FF_10;
                10'd27: pixel <= 24'hFF_12_19;
                10'd28: pixel <= 24'h09_A0_D4;
                10'd29: pixel <= 24'h66_B3_FF;
                10'd30: pixel <= 24'hAE_FF_27;
                10'd31: pixel <= 24'hFF_28_65;
                10'd32: pixel <= 24'h28_64_B0;
                10'd33: pixel <= 24'h66_B1_FF;
                10'd34: pixel <= 24'hC1_FF_29;
                10'd35: pixel <= 24'hFF_15_7E;
                10'd36: pixel <= 24'h12_1B_45;
                10'd37: pixel <= 24'h1A_42_FF;
                10'd38: pixel <= 24'h42_FF_11;
                10'd39: pixel <= 24'hFF_11_1A;
                10'd40: pixel <= 24'h0F_1B_42;
                10'd41: pixel <= 24'h1A_42_FF;
                10'd42: pixel <= 24'h44_FF_11;
                10'd43: pixel <= 24'hFF_0F_1B;
                10'd44: pixel <= 24'h1E_0E_43;
                10'd45: pixel <= 24'h2B_8A_FF;
                10'd46: pixel <= 24'hA2_FF_9C;
                10'd47: pixel <= 24'hFF_BD_5B;
                10'd48: pixel <= 24'hBD_5B_A2;
                10'd49: pixel <= 24'h5B_A2_FF;
                10'd50: pixel <= 24'hA2_FF_BB;
                10'd51: pixel <= 24'hFF_BD_5B;
                10'd52: pixel <= 24'hBC_59_A1;
                10'd53: pixel <= 24'h26_7C_FF;
                10'd54: pixel <= 24'h42_FF_84;
                10'd55: pixel <= 24'hFF_12_19;
                10'd56: pixel <= 24'h11_1A_42;
                10'd57: pixel <= 24'h1A_42_FF;
                10'd58: pixel <= 24'h42_FF_11;
                10'd59: pixel <= 24'hFF_11_1A;
                10'd60: pixel <= 24'h0E_1A_3F;
                10'd61: pixel <= 24'h4D_91_FF;
                10'd62: pixel <= 24'h8E_FF_2B;
                10'd63: pixel <= 24'hFF_24_4B;
                10'd64: pixel <= 24'h24_4A_92;
                10'd65: pixel <= 24'h41_81_FF;
                10'd66: pixel <= 24'h83_FF_22;
                10'd67: pixel <= 24'hFF_24_3F;
                10'd68: pixel <= 24'h24_49_8E;
                10'd69: pixel <= 24'h4A_8C_FF;
                10'd70: pixel <= 24'h8B_FF_23;
                10'd71: pixel <= 24'hFF_23_48;
                10'd72: pixel <= 24'h0A_1E_4C;
                10'd73: pixel <= 24'h1A_3F_FF;
                10'd74: pixel <= 24'h3F_FF_0E;
                10'd75: pixel <= 24'hFF_0E_1A;
                10'd76: pixel <= 24'h0E_1A_3F;
                10'd77: pixel <= 24'h19_3F_FF;
                10'd78: pixel <= 24'h3F_FF_10;
                10'd79: pixel <= 24'hFF_0E_1A;
                10'd80: pixel <= 24'h10_19_3F;
                10'd81: pixel <= 24'h17_3D_FF;
                10'd82: pixel <= 24'h3F_FF_14;
                10'd83: pixel <= 24'hFF_EB_25;
                10'd84: pixel <= 24'hF0_4A_65;
                10'd85: pixel <= 24'h4B_67_FF;
                10'd86: pixel <= 24'h67_FF_EF;
                10'd87: pixel <= 24'hFF_EF_4B;
                10'd88: pixel <= 24'hEF_4B_67;
                10'd89: pixel <= 24'h2A_38_FF;
                10'd90: pixel <= 24'h3F_FF_EE;
                10'd91: pixel <= 24'hFF_10_19;
                10'd92: pixel <= 24'h0E_1A_3F;
                10'd93: pixel <= 24'h1A_3F_FF;
                10'd94: pixel <= 24'h3F_FF_0E;
                10'd95: pixel <= 24'hFF_0E_1A;
                10'd96: pixel <= 24'h0D_18_42;
                10'd97: pixel <= 24'h84_1D_FF;
                10'd98: pixel <= 24'h26_FF_F0;
                10'd99: pixel <= 24'hFF_EB_30;
            endcase
            10'd7: case (x)
                10'd0: pixel <= 24'h2A_69_B3;
                10'd1: pixel <= 24'h7D_C0_FF;
                10'd2: pixel <= 24'h47_FF_14;
                10'd3: pixel <= 24'hFF_12_1D;
                10'd4: pixel <= 24'h13_1D_45;
                10'd5: pixel <= 24'h1D_45_FF;
                10'd6: pixel <= 24'h45_FF_13;
                10'd7: pixel <= 24'hFF_13_1D;
                10'd8: pixel <= 24'h13_1D_45;
                10'd9: pixel <= 24'h1D_45_FF;
                10'd10: pixel <= 24'h41_FF_13;
                10'd11: pixel <= 24'hFF_10_1D;
                10'd12: pixel <= 24'h89_42_90;
                10'd13: pixel <= 24'h2F_83_FF;
                10'd14: pixel <= 24'h58_FF_91;
                10'd15: pixel <= 24'hFF_65_17;
                10'd16: pixel <= 24'hBD_60_A6;
                10'd17: pixel <= 24'h5A_A3_FF;
                10'd18: pixel <= 24'hA3_FF_BA;
                10'd19: pixel <= 24'hFF_BA_5A;
                10'd20: pixel <= 24'hBE_59_A6;
                10'd21: pixel <= 24'h19_5D_FF;
                10'd22: pixel <= 24'h45_FF_63;
                10'd23: pixel <= 24'hFF_15_1C;
                10'd24: pixel <= 24'h15_1C_45;
                10'd25: pixel <= 24'h1D_45_FF;
                10'd26: pixel <= 24'h43_FF_13;
                10'd27: pixel <= 24'hFF_12_1E;
                10'd28: pixel <= 24'h29_4C_90;
                10'd29: pixel <= 24'h4D_92_FF;
                10'd30: pixel <= 24'h90_FF_26;
                10'd31: pixel <= 24'hFF_26_4E;
                10'd32: pixel <= 24'h22_40_83;
                10'd33: pixel <= 24'h3F_83_FF;
                10'd34: pixel <= 24'h8F_FF_24;
                10'd35: pixel <= 24'hFF_25_4C;
                10'd36: pixel <= 24'h25_4C_91;
                10'd37: pixel <= 24'h4A_8E_FF;
                10'd38: pixel <= 24'h4F_FF_26;
                10'd39: pixel <= 24'hFF_0B_1F;
                10'd40: pixel <= 24'h0F_1B_42;
                10'd41: pixel <= 24'h1A_42_FF;
                10'd42: pixel <= 24'h42_FF_11;
                10'd43: pixel <= 24'hFF_11_1A;
                10'd44: pixel <= 24'h11_1A_42;
                10'd45: pixel <= 24'h1A_42_FF;
                10'd46: pixel <= 24'h42_FF_11;
                10'd47: pixel <= 24'hFF_0F_1B;
                10'd48: pixel <= 24'h16_16_3F;
                10'd49: pixel <= 24'h25_3F_FF;
                10'd50: pixel <= 24'h67_FF_EB;
                10'd51: pixel <= 24'hFF_F0_4A;
                10'd52: pixel <= 24'hEF_4B_67;
                10'd53: pixel <= 24'h4B_67_FF;
                10'd54: pixel <= 24'h4F_FF_EF;
                10'd55: pixel <= 24'hFF_F5_3C;
                10'd56: pixel <= 24'hEE_2A_38;
                10'd57: pixel <= 24'h1A_42_FF;
                10'd58: pixel <= 24'h42_FF_11;
                10'd59: pixel <= 24'hFF_11_1A;
                10'd60: pixel <= 24'h11_1A_42;
                10'd61: pixel <= 24'h1A_42_FF;
                10'd62: pixel <= 24'h41_FF_11;
                10'd63: pixel <= 24'hFF_10_19;
                10'd64: pixel <= 24'hF0_85_21;
                10'd65: pixel <= 24'h33_24_FF;
                10'd66: pixel <= 24'h23_FF_ED;
                10'd67: pixel <= 24'hFF_EE_31;
                10'd68: pixel <= 24'hEE_31_23;
                10'd69: pixel <= 24'h33_24_FF;
                10'd70: pixel <= 24'h1E_FF_ED;
                10'd71: pixel <= 24'hFF_EE_7B;
                10'd72: pixel <= 24'h12_19_44;
                10'd73: pixel <= 24'h1A_40_FF;
                10'd74: pixel <= 24'h41_FF_12;
                10'd75: pixel <= 24'hFF_10_1D;
                10'd76: pixel <= 24'h0C_1D_3E;
                10'd77: pixel <= 24'h1A_44_FF;
                10'd78: pixel <= 24'h42_FF_11;
                10'd79: pixel <= 24'hFF_11_1A;
                10'd80: pixel <= 24'h0F_1B_42;
                10'd81: pixel <= 24'h1B_42_FF;
                10'd82: pixel <= 24'h40_FF_0F;
                10'd83: pixel <= 24'hFF_11_1B;
                10'd84: pixel <= 24'h0F_1B_42;
                10'd85: pixel <= 24'h1B_42_FF;
                10'd86: pixel <= 24'h42_FF_0F;
                10'd87: pixel <= 24'hFF_11_1A;
                10'd88: pixel <= 24'h11_1A_42;
                10'd89: pixel <= 24'h10_15_FF;
                10'd90: pixel <= 24'h21_FF_0C;
                10'd91: pixel <= 24'hFF_FF_B4;
                10'd92: pixel <= 24'hF6_8C_20;
                10'd93: pixel <= 24'h8D_1E_FF;
                10'd94: pixel <= 24'h1E_FF_F6;
                10'd95: pixel <= 24'hFF_F6_8D;
                10'd96: pixel <= 24'hF6_8D_1E;
                10'd97: pixel <= 24'hA9_41_FF;
                10'd98: pixel <= 24'h40_FF_E8;
                10'd99: pixel <= 24'hFF_11_1B;
            endcase
            10'd8: case (x)
                10'd0: pixel <= 24'h24_3F_83;
                10'd1: pixel <= 24'h4D_92_FF;
                10'd2: pixel <= 24'h92_FF_26;
                10'd3: pixel <= 24'hFF_26_4D;
                10'd4: pixel <= 24'h27_4C_8F;
                10'd5: pixel <= 24'h21_51_FF;
                10'd6: pixel <= 24'h43_FF_0D;
                10'd7: pixel <= 24'hFF_12_1B;
                10'd8: pixel <= 24'h12_1B_43;
                10'd9: pixel <= 24'h1B_43_FF;
                10'd10: pixel <= 24'h43_FF_12;
                10'd11: pixel <= 24'hFF_12_1B;
                10'd12: pixel <= 24'h12_1B_43;
                10'd13: pixel <= 24'h1B_43_FF;
                10'd14: pixel <= 24'h40_FF_12;
                10'd15: pixel <= 24'hFF_16_18;
                10'd16: pixel <= 24'hE9_24_3B;
                10'd17: pixel <= 24'h26_31_FF;
                10'd18: pixel <= 24'h27_FF_E9;
                10'd19: pixel <= 24'hFF_EE_22;
                10'd20: pixel <= 24'hEE_22_29;
                10'd21: pixel <= 24'h22_29_FF;
                10'd22: pixel <= 24'h38_FF_EE;
                10'd23: pixel <= 24'hFF_EE_2A;
                10'd24: pixel <= 24'h13_1D_45;
                10'd25: pixel <= 24'h1D_45_FF;
                10'd26: pixel <= 24'h45_FF_13;
                10'd27: pixel <= 24'hFF_13_1D;
                10'd28: pixel <= 24'h13_1D_45;
                10'd29: pixel <= 24'h1B_43_FF;
                10'd30: pixel <= 24'h1F_FF_12;
                10'd31: pixel <= 24'hFF_EF_84;
                10'd32: pixel <= 24'hEE_36_25;
                10'd33: pixel <= 24'h36_27_FF;
                10'd34: pixel <= 24'h25_FF_EE;
                10'd35: pixel <= 24'hFF_F0_35;
                10'd36: pixel <= 24'hEE_36_25;
                10'd37: pixel <= 24'h7C_1F_FF;
                10'd38: pixel <= 24'h41_FF_EF;
                10'd39: pixel <= 24'hFF_14_1B;
                10'd40: pixel <= 24'h13_1D_45;
                10'd41: pixel <= 24'h1D_45_FF;
                10'd42: pixel <= 24'h45_FF_13;
                10'd43: pixel <= 24'hFF_13_1D;
                10'd44: pixel <= 24'h13_1D_45;
                10'd45: pixel <= 24'h1D_45_FF;
                10'd46: pixel <= 24'h45_FF_13;
                10'd47: pixel <= 24'hFF_13_1D;
                10'd48: pixel <= 24'h13_1D_45;
                10'd49: pixel <= 24'h1D_45_FF;
                10'd50: pixel <= 24'h45_FF_13;
                10'd51: pixel <= 24'hFF_13_1D;
                10'd52: pixel <= 24'h13_1D_45;
                10'd53: pixel <= 24'h1D_45_FF;
                10'd54: pixel <= 24'h45_FF_13;
                10'd55: pixel <= 24'hFF_13_1D;
                10'd56: pixel <= 24'h0E_12_18;
                10'd57: pixel <= 24'hB2_24_FF;
                10'd58: pixel <= 24'h1F_FF_FF;
                10'd59: pixel <= 24'hFF_F8_8F;
                10'd60: pixel <= 24'hF8_8F_1F;
                10'd61: pixel <= 24'h8F_1F_FF;
                10'd62: pixel <= 24'h1E_FF_F8;
                10'd63: pixel <= 24'hFF_F8_8D;
                10'd64: pixel <= 24'hE8_A9_41;
                10'd65: pixel <= 24'h1D_45_FF;
                10'd66: pixel <= 24'h45_FF_13;
                10'd67: pixel <= 24'hFF_13_1D;
                10'd68: pixel <= 24'h13_1D_45;
                10'd69: pixel <= 24'h1D_45_FF;
                10'd70: pixel <= 24'h43_FF_13;
                10'd71: pixel <= 24'hFF_12_1B;
                10'd72: pixel <= 24'h52_B0_40;
                10'd73: pixel <= 24'h80_45_FF;
                10'd74: pixel <= 24'h43_FF_19;
                10'd75: pixel <= 24'hFF_18_82;
                10'd76: pixel <= 24'h19_81_43;
                10'd77: pixel <= 24'h81_41_FF;
                10'd78: pixel <= 24'h4B_FF_19;
                10'd79: pixel <= 24'hFF_48_B1;
                10'd80: pixel <= 24'h13_1C_47;
                10'd81: pixel <= 24'h1C_43_FF;
                10'd82: pixel <= 24'h49_FF_15;
                10'd83: pixel <= 24'hFF_16_1A;
                10'd84: pixel <= 24'h39_B2_50;
                10'd85: pixel <= 24'h81_41_FF;
                10'd86: pixel <= 24'h3F_FF_17;
                10'd87: pixel <= 24'hFF_18_80;
                10'd88: pixel <= 24'h18_82_43;
                10'd89: pixel <= 24'h82_41_FF;
                10'd90: pixel <= 24'h3F_FF_18;
                10'd91: pixel <= 24'hFF_18_80;
                10'd92: pixel <= 24'h21_81_38;
                10'd93: pixel <= 24'h1B_45_FF;
                10'd94: pixel <= 24'hD3_FF_12;
                10'd95: pixel <= 24'hFF_08_9F;
                10'd96: pixel <= 24'h28_69_B5;
                10'd97: pixel <= 24'h6A_B3_FF;
                10'd98: pixel <= 24'hB3_FF_28;
                10'd99: pixel <= 24'hFF_2A_69;
            endcase
            10'd9: case (x)
                10'd0: pixel <= 24'hEF_3A_25;
                10'd1: pixel <= 24'h3A_25_FF;
                10'd2: pixel <= 24'h23_FF_EF;
                10'd3: pixel <= 24'hFF_ED_3B;
                10'd4: pixel <= 24'hEC_7C_20;
                10'd5: pixel <= 24'h1D_49_FF;
                10'd6: pixel <= 24'h46_FF_12;
                10'd7: pixel <= 24'hFF_14_1E;
                10'd8: pixel <= 24'h14_1D_48;
                10'd9: pixel <= 24'h1E_46_FF;
                10'd10: pixel <= 24'h48_FF_14;
                10'd11: pixel <= 24'hFF_14_1D;
                10'd12: pixel <= 24'h14_1E_46;
                10'd13: pixel <= 24'h1D_48_FF;
                10'd14: pixel <= 24'h48_FF_14;
                10'd15: pixel <= 24'hFF_14_1D;
                10'd16: pixel <= 24'h14_1D_48;
                10'd17: pixel <= 24'h1D_48_FF;
                10'd18: pixel <= 24'h48_FF_14;
                10'd19: pixel <= 24'hFF_14_1D;
                10'd20: pixel <= 24'h14_1D_48;
                10'd21: pixel <= 24'h1D_48_FF;
                10'd22: pixel <= 24'h19_FF_14;
                10'd23: pixel <= 24'hFF_0F_13;
                10'd24: pixel <= 24'hFF_B5_21;
                10'd25: pixel <= 24'h92_1E_FF;
                10'd26: pixel <= 24'h20_FF_F8;
                10'd27: pixel <= 24'hFF_F8_91;
                10'd28: pixel <= 24'hF8_91_20;
                10'd29: pixel <= 24'h92_1F_FF;
                10'd30: pixel <= 24'h41_FF_FA;
                10'd31: pixel <= 24'hFF_E8_A9;
                10'd32: pixel <= 24'h13_1C_47;
                10'd33: pixel <= 24'h1D_48_FF;
                10'd34: pixel <= 24'h46_FF_14;
                10'd35: pixel <= 24'hFF_14_1E;
                10'd36: pixel <= 24'h14_1E_46;
                10'd37: pixel <= 24'h1E_46_FF;
                10'd38: pixel <= 24'h40_FF_14;
                10'd39: pixel <= 24'hFF_52_B0;
                10'd40: pixel <= 24'h19_85_45;
                10'd41: pixel <= 24'h86_41_FF;
                10'd42: pixel <= 24'h43_FF_17;
                10'd43: pixel <= 24'hFF_17_86;
                10'd44: pixel <= 24'h17_86_43;
                10'd45: pixel <= 24'hB3_4B_FF;
                10'd46: pixel <= 24'h46_FF_49;
                10'd47: pixel <= 24'hFF_14_1E;
                10'd48: pixel <= 24'h14_1E_44;
                10'd49: pixel <= 24'h1D_48_FF;
                10'd50: pixel <= 24'h2A_FF_14;
                10'd51: pixel <= 24'hFF_03_2F;
                10'd52: pixel <= 24'h3D_B1_51;
                10'd53: pixel <= 24'h85_43_FF;
                10'd54: pixel <= 24'h43_FF_19;
                10'd55: pixel <= 24'hFF_19_85;
                10'd56: pixel <= 24'h19_85_43;
                10'd57: pixel <= 24'h86_43_FF;
                10'd58: pixel <= 24'h3C_FF_17;
                10'd59: pixel <= 24'hFF_1E_82;
                10'd60: pixel <= 24'h15_1B_47;
                10'd61: pixel <= 24'hA2_D5_FF;
                10'd62: pixel <= 24'hB7_FF_09;
                10'd63: pixel <= 24'hFF_29_6C;
                10'd64: pixel <= 24'h28_6F_B7;
                10'd65: pixel <= 24'h6F_B7_FF;
                10'd66: pixel <= 24'hB7_FF_28;
                10'd67: pixel <= 24'hFF_28_6F;
                10'd68: pixel <= 24'h14_7D_C0;
                10'd69: pixel <= 24'h1D_48_FF;
                10'd70: pixel <= 24'h48_FF_14;
                10'd71: pixel <= 24'hFF_14_1D;
                10'd72: pixel <= 24'h14_1D_48;
                10'd73: pixel <= 24'h1E_46_FF;
                10'd74: pixel <= 24'h48_FF_14;
                10'd75: pixel <= 24'hFF_14_1D;
                10'd76: pixel <= 24'h14_1D_48;
                10'd77: pixel <= 24'h1D_48_FF;
                10'd78: pixel <= 24'h48_FF_14;
                10'd79: pixel <= 24'hFF_13_1E;
                10'd80: pixel <= 24'h98_2D_8F;
                10'd81: pixel <= 24'h21_61_FF;
                10'd82: pixel <= 24'h62_FF_6C;
                10'd83: pixel <= 24'hFF_6D_23;
                10'd84: pixel <= 24'h6D_23_62;
                10'd85: pixel <= 24'h20_61_FF;
                10'd86: pixel <= 24'hA3_FF_6F;
                10'd87: pixel <= 24'hFF_B1_5E;
                10'd88: pixel <= 24'h9B_31_8B;
                10'd89: pixel <= 24'h1B_47_FF;
                10'd90: pixel <= 24'h45_FF_15;
                10'd91: pixel <= 24'hFF_12_1D;
                10'd92: pixel <= 24'h14_1E_46;
                10'd93: pixel <= 24'h1D_43_FF;
                10'd94: pixel <= 24'h92_FF_13;
                10'd95: pixel <= 24'hFF_2C_4E;
                10'd96: pixel <= 24'h29_4F_94;
                10'd97: pixel <= 24'h51_92_FF;
                10'd98: pixel <= 24'h83_FF_27;
                10'd99: pixel <= 24'hFF_22_40;
            endcase
            10'd10: case (x)
                10'd0: pixel <= 24'h17_1E_49;
                10'd1: pixel <= 24'h1E_49_FF;
                10'd2: pixel <= 24'h49_FF_17;
                10'd3: pixel <= 24'hFF_17_1E;
                10'd4: pixel <= 24'h17_1E_49;
                10'd5: pixel <= 24'hAF_40_FF;
                10'd6: pixel <= 24'h44_FF_54;
                10'd7: pixel <= 24'hFF_18_87;
                10'd8: pixel <= 24'h18_88_42;
                10'd9: pixel <= 24'h88_42_FF;
                10'd10: pixel <= 24'h46_FF_18;
                10'd11: pixel <= 24'hFF_18_87;
                10'd12: pixel <= 24'h48_B1_49;
                10'd13: pixel <= 24'h20_48_FF;
                10'd14: pixel <= 24'h47_FF_17;
                10'd15: pixel <= 24'hFF_17_1E;
                10'd16: pixel <= 24'h15_1E_49;
                10'd17: pixel <= 24'h1F_48_FF;
                10'd18: pixel <= 24'h4D_FF_18;
                10'd19: pixel <= 24'hFF_35_A2;
                10'd20: pixel <= 24'h1A_8B_3B;
                10'd21: pixel <= 24'h88_42_FF;
                10'd22: pixel <= 24'h42_FF_18;
                10'd23: pixel <= 24'hFF_18_88;
                10'd24: pixel <= 24'h18_88_42;
                10'd25: pixel <= 24'h82_3A_FF;
                10'd26: pixel <= 24'h48_FF_1E;
                10'd27: pixel <= 24'hFF_16_1C;
                10'd28: pixel <= 24'h09_A2_D5;
                10'd29: pixel <= 24'h6F_BA_FF;
                10'd30: pixel <= 24'hB8_FF_2A;
                10'd31: pixel <= 24'hFF_28_71;
                10'd32: pixel <= 24'h28_71_B8;
                10'd33: pixel <= 24'h72_B9_FF;
                10'd34: pixel <= 24'hC0_FF_29;
                10'd35: pixel <= 24'hFF_12_7E;
                10'd36: pixel <= 24'h15_1E_49;
                10'd37: pixel <= 24'h55_A0_FF;
                10'd38: pixel <= 24'hA1_FF_B8;
                10'd39: pixel <= 24'hFF_B4_4F;
                10'd40: pixel <= 24'hAF_48_9D;
                10'd41: pixel <= 24'h43_9B_FF;
                10'd42: pixel <= 24'h9B_FF_AB;
                10'd43: pixel <= 24'hFF_A8_3F;
                10'd44: pixel <= 24'hA4_39_97;
                10'd45: pixel <= 24'h33_94_FF;
                10'd46: pixel <= 24'h85_FF_A1;
                10'd47: pixel <= 24'hFF_8C_2F;
                10'd48: pixel <= 24'h6E_21_64;
                10'd49: pixel <= 24'h21_64_FF;
                10'd50: pixel <= 24'h64_FF_6E;
                10'd51: pixel <= 24'hFF_6E_21;
                10'd52: pixel <= 24'h6E_21_64;
                10'd53: pixel <= 24'h21_60_FF;
                10'd54: pixel <= 24'h8C_FF_70;
                10'd55: pixel <= 24'hFF_9B_2F;
                10'd56: pixel <= 24'h1B_1A_48;
                10'd57: pixel <= 24'h1D_48_FF;
                10'd58: pixel <= 24'h48_FF_14;
                10'd59: pixel <= 24'hFF_16_1C;
                10'd60: pixel <= 24'h15_1C_45;
                10'd61: pixel <= 24'h4E_91_FF;
                10'd62: pixel <= 24'h95_FF_29;
                10'd63: pixel <= 24'hFF_2A_51;
                10'd64: pixel <= 24'h2A_50_99;
                10'd65: pixel <= 24'h40_83_FF;
                10'd66: pixel <= 24'h83_FF_22;
                10'd67: pixel <= 24'hFF_24_3F;
                10'd68: pixel <= 24'h29_4F_94;
                10'd69: pixel <= 24'h4F_94_FF;
                10'd70: pixel <= 24'h93_FF_29;
                10'd71: pixel <= 24'hFF_2B_50;
                10'd72: pixel <= 24'h10_23_53;
                10'd73: pixel <= 24'h1E_46_FF;
                10'd74: pixel <= 24'h48_FF_14;
                10'd75: pixel <= 24'hFF_14_1D;
                10'd76: pixel <= 24'h14_1D_48;
                10'd77: pixel <= 24'h1D_48_FF;
                10'd78: pixel <= 24'h46_FF_14;
                10'd79: pixel <= 24'hFF_14_1E;
                10'd80: pixel <= 24'h14_1E_46;
                10'd81: pixel <= 24'h1A_3F_FF;
                10'd82: pixel <= 24'h35_FF_17;
                10'd83: pixel <= 24'hFF_EE_23;
                10'd84: pixel <= 24'hEF_23_28;
                10'd85: pixel <= 24'h22_27_FF;
                10'd86: pixel <= 24'h27_FF_EE;
                10'd87: pixel <= 24'hFF_EE_22;
                10'd88: pixel <= 24'hEF_21_29;
                10'd89: pixel <= 24'h2A_38_FF;
                10'd90: pixel <= 24'h46_FF_EE;
                10'd91: pixel <= 24'hFF_14_1E;
                10'd92: pixel <= 24'h14_1D_48;
                10'd93: pixel <= 24'h1D_48_FF;
                10'd94: pixel <= 24'h48_FF_14;
                10'd95: pixel <= 24'hFF_14_1D;
                10'd96: pixel <= 24'h13_1C_47;
                10'd97: pixel <= 24'h83_1E_FF;
                10'd98: pixel <= 24'h22_FF_EE;
                10'd99: pixel <= 24'hFF_EC_3A;
            endcase
            10'd11: case (x)
                10'd0: pixel <= 24'h25_75_BA;
                10'd1: pixel <= 24'h7E_C0_FF;
                10'd2: pixel <= 24'h4D_FF_12;
                10'd3: pixel <= 24'hFF_19_20;
                10'd4: pixel <= 24'hB8_50_A0;
                10'd5: pixel <= 24'h23_69_FF;
                10'd6: pixel <= 24'h67_FF_72;
                10'd7: pixel <= 24'hFF_72_23;
                10'd8: pixel <= 24'h74_22_69;
                10'd9: pixel <= 24'h21_6B_FF;
                10'd10: pixel <= 24'h69_FF_74;
                10'd11: pixel <= 24'hFF_72_23;
                10'd12: pixel <= 24'h72_23_69;
                10'd13: pixel <= 24'h23_69_FF;
                10'd14: pixel <= 24'h69_FF_72;
                10'd15: pixel <= 24'hFF_71_23;
                10'd16: pixel <= 24'h72_23_67;
                10'd17: pixel <= 24'h23_69_FF;
                10'd18: pixel <= 24'h69_FF_72;
                10'd19: pixel <= 24'hFF_72_23;
                10'd20: pixel <= 24'h72_22_6D;
                10'd21: pixel <= 24'h2D_8E_FF;
                10'd22: pixel <= 24'h4B_FF_9D;
                10'd23: pixel <= 24'hFF_19_1C;
                10'd24: pixel <= 24'h18_1F_4A;
                10'd25: pixel <= 24'h1F_4A_FF;
                10'd26: pixel <= 24'h49_FF_18;
                10'd27: pixel <= 24'hFF_16_22;
                10'd28: pixel <= 24'h2F_51_98;
                10'd29: pixel <= 24'h51_99_FF;
                10'd30: pixel <= 24'h9B_FF_2B;
                10'd31: pixel <= 24'hFF_29_52;
                10'd32: pixel <= 24'h22_40_83;
                10'd33: pixel <= 24'h3F_83_FF;
                10'd34: pixel <= 24'h94_FF_24;
                10'd35: pixel <= 24'hFF_29_4F;
                10'd36: pixel <= 24'h2A_51_95;
                10'd37: pixel <= 24'h50_93_FF;
                10'd38: pixel <= 24'h53_FF_2B;
                10'd39: pixel <= 24'hFF_10_23;
                10'd40: pixel <= 24'h14_1D_48;
                10'd41: pixel <= 24'h1C_48_FF;
                10'd42: pixel <= 24'h49_FF_16;
                10'd43: pixel <= 24'hFF_17_1E;
                10'd44: pixel <= 24'h17_1E_49;
                10'd45: pixel <= 24'h1E_49_FF;
                10'd46: pixel <= 24'h49_FF_17;
                10'd47: pixel <= 24'hFF_17_1E;
                10'd48: pixel <= 24'h1A_1D_45;
                10'd49: pixel <= 24'h24_37_FF;
                10'd50: pixel <= 24'h27_FF_EF;
                10'd51: pixel <= 24'hFF_EE_22;
                10'd52: pixel <= 24'hEE_22_27;
                10'd53: pixel <= 24'h22_27_FF;
                10'd54: pixel <= 24'h29_FF_EE;
                10'd55: pixel <= 24'hFF_EF_21;
                10'd56: pixel <= 24'hEE_2A_38;
                10'd57: pixel <= 24'h1E_49_FF;
                10'd58: pixel <= 24'h49_FF_17;
                10'd59: pixel <= 24'hFF_17_1E;
                10'd60: pixel <= 24'h17_1E_49;
                10'd61: pixel <= 24'h1E_49_FF;
                10'd62: pixel <= 24'h48_FF_17;
                10'd63: pixel <= 24'hFF_16_1C;
                10'd64: pixel <= 24'hEF_84_1F;
                10'd65: pixel <= 24'h3C_24_FF;
                10'd66: pixel <= 24'h22_FF_EE;
                10'd67: pixel <= 24'hFF_ED_3D;
                10'd68: pixel <= 24'hED_3D_22;
                10'd69: pixel <= 24'h3E_20_FF;
                10'd70: pixel <= 24'h2D_FF_EB;
                10'd71: pixel <= 24'hFF_F8_62;
                10'd72: pixel <= 24'hFB_90_2D;
                10'd73: pixel <= 24'h89_25_FF;
                10'd74: pixel <= 24'h23_FF_F9;
                10'd75: pixel <= 24'hFF_F9_7F;
                10'd76: pixel <= 24'hF2_78_21;
                10'd77: pixel <= 24'h71_22_FF;
                10'd78: pixel <= 24'h1E_FF_F1;
                10'd79: pixel <= 24'hFF_EE_6A;
                10'd80: pixel <= 24'hF0_5F_21;
                10'd81: pixel <= 24'h57_21_FF;
                10'd82: pixel <= 24'h21_FF_F0;
                10'd83: pixel <= 24'hFF_ED_53;
                10'd84: pixel <= 24'h1E_19_41;
                10'd85: pixel <= 24'h1C_48_FF;
                10'd86: pixel <= 24'h48_FF_16;
                10'd87: pixel <= 24'hFF_16_1C;
                10'd88: pixel <= 24'h15_1E_49;
                10'd89: pixel <= 24'h15_1D_FF;
                10'd90: pixel <= 24'h20_FF_12;
                10'd91: pixel <= 24'hFF_FF_B3;
                10'd92: pixel <= 24'hF7_94_1D;
                10'd93: pixel <= 24'h94_1F_FF;
                10'd94: pixel <= 24'h1D_FF_F7;
                10'd95: pixel <= 24'hFF_F7_94;
                10'd96: pixel <= 24'hFA_94_20;
                10'd97: pixel <= 24'hA9_41_FF;
                10'd98: pixel <= 24'h49_FF_E8;
                10'd99: pixel <= 24'hFF_15_1E;
            endcase
            10'd12: case (x)
                10'd0: pixel <= 24'h24_3F_83;
                10'd1: pixel <= 24'h51_99_FF;
                10'd2: pixel <= 24'h9A_FF_2B;
                10'd3: pixel <= 24'hFF_2C_53;
                10'd4: pixel <= 24'h2F_51_98;
                10'd5: pixel <= 24'h23_57_FF;
                10'd6: pixel <= 24'h4A_FF_13;
                10'd7: pixel <= 24'hFF_18_1F;
                10'd8: pixel <= 24'h18_1E_4C;
                10'd9: pixel <= 24'h1E_4C_FF;
                10'd10: pixel <= 24'h4C_FF_18;
                10'd11: pixel <= 24'hFF_18_1E;
                10'd12: pixel <= 24'h18_1F_4A;
                10'd13: pixel <= 24'h1E_4C_FF;
                10'd14: pixel <= 24'h47_FF_18;
                10'd15: pixel <= 24'hFF_1A_1C;
                10'd16: pixel <= 24'hEF_24_35;
                10'd17: pixel <= 24'h22_27_FF;
                10'd18: pixel <= 24'h27_FF_EE;
                10'd19: pixel <= 24'hFF_EE_22;
                10'd20: pixel <= 24'hEE_22_27;
                10'd21: pixel <= 24'h20_2B_FF;
                10'd22: pixel <= 24'h38_FF_EF;
                10'd23: pixel <= 24'hFF_EE_2A;
                10'd24: pixel <= 24'h18_1E_4C;
                10'd25: pixel <= 24'h1F_4A_FF;
                10'd26: pixel <= 24'h4A_FF_18;
                10'd27: pixel <= 24'hFF_18_1F;
                10'd28: pixel <= 24'h18_1E_4C;
                10'd29: pixel <= 24'h1E_49_FF;
                10'd30: pixel <= 24'h1E_FF_17;
                10'd31: pixel <= 24'hFF_F0_8C;
                10'd32: pixel <= 24'hED_40_24;
                10'd33: pixel <= 24'h41_22_FF;
                10'd34: pixel <= 24'h24_FF_ED;
                10'd35: pixel <= 24'hFF_ED_40;
                10'd36: pixel <= 24'hED_40_24;
                10'd37: pixel <= 24'h41_22_FF;
                10'd38: pixel <= 24'h21_FF_ED;
                10'd39: pixel <= 24'hFF_EC_40;
                10'd40: pixel <= 24'hED_40_24;
                10'd41: pixel <= 24'h40_24_FF;
                10'd42: pixel <= 24'h24_FF_ED;
                10'd43: pixel <= 24'hFF_ED_40;
                10'd44: pixel <= 24'hED_40_24;
                10'd45: pixel <= 24'h40_24_FF;
                10'd46: pixel <= 24'h24_FF_ED;
                10'd47: pixel <= 24'hFF_ED_40;
                10'd48: pixel <= 24'hED_41_22;
                10'd49: pixel <= 24'h44_1F_FF;
                10'd50: pixel <= 24'h28_FF_F0;
                10'd51: pixel <= 24'hFF_E7_4B;
                10'd52: pixel <= 24'h1B_1D_4A;
                10'd53: pixel <= 24'h1D_49_FF;
                10'd54: pixel <= 24'h4A_FF_19;
                10'd55: pixel <= 24'hFF_18_1F;
                10'd56: pixel <= 24'h15_15_20;
                10'd57: pixel <= 24'hB4_1F_FF;
                10'd58: pixel <= 24'h1D_FF_FB;
                10'd59: pixel <= 24'hFF_F6_98;
                10'd60: pixel <= 24'hF8_98_1D;
                10'd61: pixel <= 24'h98_1D_FF;
                10'd62: pixel <= 24'h1D_FF_F6;
                10'd63: pixel <= 24'hFF_F8_98;
                10'd64: pixel <= 24'hE8_A9_3F;
                10'd65: pixel <= 24'h1E_4C_FF;
                10'd66: pixel <= 24'h4A_FF_18;
                10'd67: pixel <= 24'hFF_18_1F;
                10'd68: pixel <= 24'h18_1E_4C;
                10'd69: pixel <= 24'h1E_4C_FF;
                10'd70: pixel <= 24'h4C_FF_18;
                10'd71: pixel <= 24'hFF_18_1E;
                10'd72: pixel <= 24'h54_AE_44;
                10'd73: pixel <= 24'h8B_44_FF;
                10'd74: pixel <= 24'h42_FF_19;
                10'd75: pixel <= 24'hFF_19_8B;
                10'd76: pixel <= 24'h19_8B_44;
                10'd77: pixel <= 24'h8B_44_FF;
                10'd78: pixel <= 24'h4B_FF_19;
                10'd79: pixel <= 24'hFF_48_B1;
                10'd80: pixel <= 24'h17_20_4A;
                10'd81: pixel <= 24'h1F_4A_FF;
                10'd82: pixel <= 24'h4A_FF_18;
                10'd83: pixel <= 24'hFF_18_1F;
                10'd84: pixel <= 24'h18_1F_4A;
                10'd85: pixel <= 24'h23_43_FF;
                10'd86: pixel <= 24'h4E_FF_13;
                10'd87: pixel <= 24'hFF_3E_B0;
                10'd88: pixel <= 24'h19_8B_40;
                10'd89: pixel <= 24'h8B_42_FF;
                10'd90: pixel <= 24'h44_FF_19;
                10'd91: pixel <= 24'hFF_19_8B;
                10'd92: pixel <= 24'h1C_83_3A;
                10'd93: pixel <= 24'h20_48_FF;
                10'd94: pixel <= 24'hD2_FF_17;
                10'd95: pixel <= 24'hFF_05_9F;
                10'd96: pixel <= 24'h24_76_BC;
                10'd97: pixel <= 24'h75_BC_FF;
                10'd98: pixel <= 24'hBA_FF_25;
                10'd99: pixel <= 24'hFF_25_75;
            endcase
            10'd13: case (x)
                10'd0: pixel <= 24'hEE_44_23;
                10'd1: pixel <= 24'h44_25_FF;
                10'd2: pixel <= 24'h23_FF_EE;
                10'd3: pixel <= 24'hFF_EE_44;
                10'd4: pixel <= 24'hEE_44_23;
                10'd5: pixel <= 24'h44_23_FF;
                10'd6: pixel <= 24'h24_FF_EE;
                10'd7: pixel <= 24'hFF_EE_46;
                10'd8: pixel <= 24'hEF_46_24;
                10'd9: pixel <= 24'h46_24_FF;
                10'd10: pixel <= 24'h24_FF_EF;
                10'd11: pixel <= 24'hFF_EF_46;
                10'd12: pixel <= 24'hEF_46_24;
                10'd13: pixel <= 24'h46_24_FF;
                10'd14: pixel <= 24'h24_FF_EF;
                10'd15: pixel <= 24'hFF_EF_46;
                10'd16: pixel <= 24'hEE_44_23;
                10'd17: pixel <= 24'h6D_25_FF;
                10'd18: pixel <= 24'h34_FF_F4;
                10'd19: pixel <= 24'hFF_45_18;
                10'd20: pixel <= 24'h19_20_4B;
                10'd21: pixel <= 24'h1F_4D_FF;
                10'd22: pixel <= 24'h25_FF_1B;
                10'd23: pixel <= 24'hFF_17_17;
                10'd24: pixel <= 24'hFF_B6_1F;
                10'd25: pixel <= 24'h9C_1E_FF;
                10'd26: pixel <= 24'h1E_FF_F7;
                10'd27: pixel <= 24'hFF_F9_9B;
                10'd28: pixel <= 24'hF7_9C_1C;
                10'd29: pixel <= 24'h9A_1C_FF;
                10'd30: pixel <= 24'h3F_FF_F7;
                10'd31: pixel <= 24'hFF_E8_A9;
                10'd32: pixel <= 24'h1B_1E_4F;
                10'd33: pixel <= 24'h20_4D_FF;
                10'd34: pixel <= 24'h4D_FF_19;
                10'd35: pixel <= 24'hFF_19_20;
                10'd36: pixel <= 24'h19_20_4D;
                10'd37: pixel <= 24'h20_4D_FF;
                10'd38: pixel <= 24'h44_FF_19;
                10'd39: pixel <= 24'hFF_54_AE;
                10'd40: pixel <= 24'h1A_8E_45;
                10'd41: pixel <= 24'h8F_45_FF;
                10'd42: pixel <= 24'h43_FF_18;
                10'd43: pixel <= 24'hFF_18_8F;
                10'd44: pixel <= 24'h16_90_45;
                10'd45: pixel <= 24'hB1_4D_FF;
                10'd46: pixel <= 24'h4B_FF_48;
                10'd47: pixel <= 24'hFF_18_21;
                10'd48: pixel <= 24'h19_20_4B;
                10'd49: pixel <= 24'h20_4D_FF;
                10'd50: pixel <= 24'h4D_FF_19;
                10'd51: pixel <= 24'hFF_19_20;
                10'd52: pixel <= 24'h1B_1F_4B;
                10'd53: pixel <= 24'h8B_5E_FF;
                10'd54: pixel <= 24'h50_FF_3D;
                10'd55: pixel <= 24'hFF_33_A4;
                10'd56: pixel <= 24'h1A_8E_45;
                10'd57: pixel <= 24'h8F_45_FF;
                10'd58: pixel <= 24'h3A_FF_18;
                10'd59: pixel <= 24'hFF_1B_84;
                10'd60: pixel <= 24'h19_20_4B;
                10'd61: pixel <= 24'hA1_D4_FF;
                10'd62: pixel <= 24'hBF_FF_08;
                10'd63: pixel <= 24'hFF_23_77;
                10'd64: pixel <= 24'h26_78_BE;
                10'd65: pixel <= 24'h77_BE_FF;
                10'd66: pixel <= 24'hBB_FF_28;
                10'd67: pixel <= 24'hFF_27_77;
                10'd68: pixel <= 24'h12_7E_C0;
                10'd69: pixel <= 24'h1F_4F_FF;
                10'd70: pixel <= 24'hA0_FF_19;
                10'd71: pixel <= 24'hFF_B8_50;
                10'd72: pixel <= 24'h76_24_6B;
                10'd73: pixel <= 24'h24_6D_FF;
                10'd74: pixel <= 24'h6D_FF_76;
                10'd75: pixel <= 24'hFF_76_24;
                10'd76: pixel <= 24'h76_24_6D;
                10'd77: pixel <= 24'h24_6D_FF;
                10'd78: pixel <= 24'h6D_FF_76;
                10'd79: pixel <= 24'hFF_76_24;
                10'd80: pixel <= 24'h76_24_6D;
                10'd81: pixel <= 24'h24_6D_FF;
                10'd82: pixel <= 24'h6D_FF_76;
                10'd83: pixel <= 24'hFF_76_24;
                10'd84: pixel <= 24'h76_24_6D;
                10'd85: pixel <= 24'h24_6D_FF;
                10'd86: pixel <= 24'h6B_FF_76;
                10'd87: pixel <= 24'hFF_76_24;
                10'd88: pixel <= 24'h8C_28_81;
                10'd89: pixel <= 24'h1F_4E_FF;
                10'd90: pixel <= 24'h4D_FF_17;
                10'd91: pixel <= 24'hFF_19_20;
                10'd92: pixel <= 24'h19_20_4D;
                10'd93: pixel <= 24'h21_49_FF;
                10'd94: pixel <= 24'h99_FF_18;
                10'd95: pixel <= 24'hFF_30_52;
                10'd96: pixel <= 24'h2C_53_9A;
                10'd97: pixel <= 24'h55_9B_FF;
                10'd98: pixel <= 24'h81_FF_2C;
                10'd99: pixel <= 24'hFF_22_41;
            endcase
            10'd14: case (x)
                10'd0: pixel <= 24'h1C_22_50;
                10'd1: pixel <= 24'h22_50_FF;
                10'd2: pixel <= 24'h50_FF_1C;
                10'd3: pixel <= 24'hFF_1C_22;
                10'd4: pixel <= 24'h1C_22_50;
                10'd5: pixel <= 24'hAE_44_FF;
                10'd6: pixel <= 24'h45_FF_54;
                10'd7: pixel <= 24'hFF_19_93;
                10'd8: pixel <= 24'h19_93_45;
                10'd9: pixel <= 24'h93_45_FF;
                10'd10: pixel <= 24'h47_FF_19;
                10'd11: pixel <= 24'hFF_19_92;
                10'd12: pixel <= 24'h48_B1_4B;
                10'd13: pixel <= 24'h23_4E_FF;
                10'd14: pixel <= 24'h4E_FF_1A;
                10'd15: pixel <= 24'hFF_1D_21;
                10'd16: pixel <= 24'h1C_22_50;
                10'd17: pixel <= 24'h22_50_FF;
                10'd18: pixel <= 24'h50_FF_1C;
                10'd19: pixel <= 24'hFF_1C_22;
                10'd20: pixel <= 24'h1D_21_50;
                10'd21: pixel <= 24'h99_40_FF;
                10'd22: pixel <= 24'h45_FF_2B;
                10'd23: pixel <= 24'hFF_18_91;
                10'd24: pixel <= 24'h18_91_46;
                10'd25: pixel <= 24'h83_38_FF;
                10'd26: pixel <= 24'h4E_FF_1E;
                10'd27: pixel <= 24'hFF_1C_20;
                10'd28: pixel <= 24'h09_A2_D7;
                10'd29: pixel <= 24'h7B_C2_FF;
                10'd30: pixel <= 24'hC1_FF_24;
                10'd31: pixel <= 24'hFF_24_7D;
                10'd32: pixel <= 24'h24_7D_C1;
                10'd33: pixel <= 24'h7C_C0_FF;
                10'd34: pixel <= 24'hC2_FF_23;
                10'd35: pixel <= 24'hFF_11_7E;
                10'd36: pixel <= 24'h1C_22_50;
                10'd37: pixel <= 24'h50_9E_FF;
                10'd38: pixel <= 24'h6E_FF_B8;
                10'd39: pixel <= 24'hFF_79_24;
                10'd40: pixel <= 24'h7A_25_71;
                10'd41: pixel <= 24'h26_71_FF;
                10'd42: pixel <= 24'h71_FF_79;
                10'd43: pixel <= 24'hFF_79_26;
                10'd44: pixel <= 24'h7A_25_71;
                10'd45: pixel <= 24'h25_71_FF;
                10'd46: pixel <= 24'h71_FF_7A;
                10'd47: pixel <= 24'hFF_7A_25;
                10'd48: pixel <= 24'h79_26_71;
                10'd49: pixel <= 24'h26_71_FF;
                10'd50: pixel <= 24'h71_FF_79;
                10'd51: pixel <= 24'hFF_7A_25;
                10'd52: pixel <= 24'h7A_25_6F;
                10'd53: pixel <= 24'h29_82_FF;
                10'd54: pixel <= 24'h5D_FF_94;
                10'd55: pixel <= 24'hFF_5B_1F;
                10'd56: pixel <= 24'h1B_21_4E;
                10'd57: pixel <= 24'h21_4E_FF;
                10'd58: pixel <= 24'h4E_FF_1B;
                10'd59: pixel <= 24'hFF_1B_21;
                10'd60: pixel <= 24'h19_22_4A;
                10'd61: pixel <= 24'h54_9A_FF;
                10'd62: pixel <= 24'h9C_FF_32;
                10'd63: pixel <= 24'hFF_2D_56;
                10'd64: pixel <= 24'h2D_56_9C;
                10'd65: pixel <= 24'h41_81_FF;
                10'd66: pixel <= 24'h81_FF_22;
                10'd67: pixel <= 24'hFF_24_40;
                10'd68: pixel <= 24'h2C_53_9A;
                10'd69: pixel <= 24'h53_9A_FF;
                10'd70: pixel <= 24'h99_FF_2C;
                10'd71: pixel <= 24'hFF_30_52;
                10'd72: pixel <= 24'h14_24_58;
                10'd73: pixel <= 24'h20_4D_FF;
                10'd74: pixel <= 24'h4D_FF_19;
                10'd75: pixel <= 24'hFF_19_20;
                10'd76: pixel <= 24'h19_20_4D;
                10'd77: pixel <= 24'h20_4D_FF;
                10'd78: pixel <= 24'h4D_FF_19;
                10'd79: pixel <= 24'hFF_19_20;
                10'd80: pixel <= 24'h19_20_4D;
                10'd81: pixel <= 24'h1C_49_FF;
                10'd82: pixel <= 24'h35_FF_1A;
                10'd83: pixel <= 24'hFF_EF_24;
                10'd84: pixel <= 24'hEE_22_27;
                10'd85: pixel <= 24'h22_27_FF;
                10'd86: pixel <= 24'h27_FF_EE;
                10'd87: pixel <= 24'hFF_EE_22;
                10'd88: pixel <= 24'hEF_23_2A;
                10'd89: pixel <= 24'h2A_3A_FF;
                10'd90: pixel <= 24'h4D_FF_EE;
                10'd91: pixel <= 24'hFF_19_20;
                10'd92: pixel <= 24'h19_20_4D;
                10'd93: pixel <= 24'h20_4D_FF;
                10'd94: pixel <= 24'h4D_FF_19;
                10'd95: pixel <= 24'hFF_19_20;
                10'd96: pixel <= 24'h19_20_4D;
                10'd97: pixel <= 24'hCC_32_FF;
                10'd98: pixel <= 24'h23_FF_FF;
                10'd99: pixel <= 24'hFF_ED_43;
            endcase
            10'd15: case (x)
                10'd0: pixel <= 24'h21_7E_C4;
                10'd1: pixel <= 24'h7F_C3_FF;
                10'd2: pixel <= 24'h50_FF_12;
                10'd3: pixel <= 24'hFF_1C_22;
                10'd4: pixel <= 24'hB8_50_A0;
                10'd5: pixel <= 24'h27_74_FF;
                10'd6: pixel <= 24'h74_FF_7A;
                10'd7: pixel <= 24'hFF_7C_26;
                10'd8: pixel <= 24'h7C_26_75;
                10'd9: pixel <= 24'h26_75_FF;
                10'd10: pixel <= 24'h75_FF_7C;
                10'd11: pixel <= 24'hFF_7C_26;
                10'd12: pixel <= 24'h7C_26_75;
                10'd13: pixel <= 24'h26_75_FF;
                10'd14: pixel <= 24'h75_FF_7C;
                10'd15: pixel <= 24'hFF_7A_26;
                10'd16: pixel <= 24'h7A_26_75;
                10'd17: pixel <= 24'h25_71_FF;
                10'd18: pixel <= 24'h85_FF_7A;
                10'd19: pixel <= 24'hFF_92_28;
                10'd20: pixel <= 24'h69_1D_62;
                10'd21: pixel <= 24'h23_52_FF;
                10'd22: pixel <= 24'h51_FF_1D;
                10'd23: pixel <= 24'hFF_1F_21;
                10'd24: pixel <= 24'h1C_22_51;
                10'd25: pixel <= 24'h22_51_FF;
                10'd26: pixel <= 24'h4C_FF_1C;
                10'd27: pixel <= 24'hFF_19_22;
                10'd28: pixel <= 24'h32_57_9C;
                10'd29: pixel <= 24'h57_9D_FF;
                10'd30: pixel <= 24'h9B_FF_2E;
                10'd31: pixel <= 24'hFF_2E_57;
                10'd32: pixel <= 24'h22_41_81;
                10'd33: pixel <= 24'h40_81_FF;
                10'd34: pixel <= 24'h9C_FF_24;
                10'd35: pixel <= 24'hFF_2D_56;
                10'd36: pixel <= 24'h2E_55_9C;
                10'd37: pixel <= 24'h53_99_FF;
                10'd38: pixel <= 24'h5B_FF_2F;
                10'd39: pixel <= 24'hFF_16_29;
                10'd40: pixel <= 24'h1B_21_4E;
                10'd41: pixel <= 24'h21_4E_FF;
                10'd42: pixel <= 24'h4E_FF_1B;
                10'd43: pixel <= 24'hFF_1B_21;
                10'd44: pixel <= 24'h1B_21_4E;
                10'd45: pixel <= 24'h22_50_FF;
                10'd46: pixel <= 24'h50_FF_1C;
                10'd47: pixel <= 24'hFF_1C_22;
                10'd48: pixel <= 24'h1E_20_4C;
                10'd49: pixel <= 24'h23_33_FF;
                10'd50: pixel <= 24'h27_FF_EE;
                10'd51: pixel <= 24'hFF_EE_22;
                10'd52: pixel <= 24'hEE_22_27;
                10'd53: pixel <= 24'h22_27_FF;
                10'd54: pixel <= 24'h2A_FF_EE;
                10'd55: pixel <= 24'hFF_EF_23;
                10'd56: pixel <= 24'hEE_2A_3A;
                10'd57: pixel <= 24'h22_50_FF;
                10'd58: pixel <= 24'h50_FF_1C;
                10'd59: pixel <= 24'hFF_1C_22;
                10'd60: pixel <= 24'h1C_22_50;
                10'd61: pixel <= 24'h22_50_FF;
                10'd62: pixel <= 24'h50_FF_1C;
                10'd63: pixel <= 24'hFF_1C_22;
                10'd64: pixel <= 24'h59_48_1F;
                10'd65: pixel <= 24'h70_29_FF;
                10'd66: pixel <= 24'h25_FF_F9;
                10'd67: pixel <= 24'hFF_EF_47;
                10'd68: pixel <= 24'hED_49_23;
                10'd69: pixel <= 24'h48_23_FF;
                10'd70: pixel <= 24'h23_FF_EF;
                10'd71: pixel <= 24'hFF_EF_48;
                10'd72: pixel <= 24'hEF_48_23;
                10'd73: pixel <= 24'h4A_24_FF;
                10'd74: pixel <= 24'h24_FF_EE;
                10'd75: pixel <= 24'hFF_F0_49;
                10'd76: pixel <= 24'hF0_49_24;
                10'd77: pixel <= 24'h49_24_FF;
                10'd78: pixel <= 24'h24_FF_F0;
                10'd79: pixel <= 24'hFF_F0_49;
                10'd80: pixel <= 24'hF0_49_24;
                10'd81: pixel <= 24'h4A_24_FF;
                10'd82: pixel <= 24'h23_FF_EE;
                10'd83: pixel <= 24'hFF_ED_49;
                10'd84: pixel <= 24'hED_49_23;
                10'd85: pixel <= 24'h47_1D_FF;
                10'd86: pixel <= 24'h4D_FF_E6;
                10'd87: pixel <= 24'hFF_1A_1E;
                10'd88: pixel <= 24'h1C_22_52;
                10'd89: pixel <= 24'h17_25_FF;
                10'd90: pixel <= 24'h1D_FF_17;
                10'd91: pixel <= 24'hFF_FD_B3;
                10'd92: pixel <= 24'hF9_9F_1C;
                10'd93: pixel <= 24'h9F_1E_FF;
                10'd94: pixel <= 24'h1E_FF_F9;
                10'd95: pixel <= 24'hFF_F8_A0;
                10'd96: pixel <= 24'hF9_9F_1E;
                10'd97: pixel <= 24'hA9_3F_FF;
                10'd98: pixel <= 24'h52_FF_E8;
                10'd99: pixel <= 24'hFF_1C_22;
            endcase
            10'd16: case (x)
                10'd0: pixel <= 24'h22_41_81;
                10'd1: pixel <= 24'h57_9D_FF;
                10'd2: pixel <= 24'h9D_FF_2E;
                10'd3: pixel <= 24'hFF_30_57;
                10'd4: pixel <= 24'h32_57_9D;
                10'd5: pixel <= 24'h28_5B_FF;
                10'd6: pixel <= 24'h50_FF_17;
                10'd7: pixel <= 24'hFF_1C_22;
                10'd8: pixel <= 24'h1C_22_51;
                10'd9: pixel <= 24'h22_51_FF;
                10'd10: pixel <= 24'h51_FF_1C;
                10'd11: pixel <= 24'hFF_1D_22;
                10'd12: pixel <= 24'h1D_23_52;
                10'd13: pixel <= 24'h23_52_FF;
                10'd14: pixel <= 24'h4B_FF_1D;
                10'd15: pixel <= 24'hFF_1D_1E;
                10'd16: pixel <= 24'hEF_24_35;
                10'd17: pixel <= 24'h22_27_FF;
                10'd18: pixel <= 24'h27_FF_EE;
                10'd19: pixel <= 24'hFF_EE_22;
                10'd20: pixel <= 24'hEC_23_27;
                10'd21: pixel <= 24'h22_2B_FF;
                10'd22: pixel <= 24'h38_FF_EF;
                10'd23: pixel <= 24'hFF_EE_2A;
                10'd24: pixel <= 24'h1D_22_51;
                10'd25: pixel <= 24'h22_51_FF;
                10'd26: pixel <= 24'h51_FF_1C;
                10'd27: pixel <= 24'hFF_1C_22;
                10'd28: pixel <= 24'h1C_22_51;
                10'd29: pixel <= 24'h22_51_FF;
                10'd30: pixel <= 24'h54_FF_1D;
                10'd31: pixel <= 24'hFF_1D_25;
                10'd32: pixel <= 24'hF3_C6_43;
                10'd33: pixel <= 24'h6A_29_FF;
                10'd34: pixel <= 24'h25_FF_F9;
                10'd35: pixel <= 24'hFF_ED_4B;
                10'd36: pixel <= 24'hEE_4A_23;
                10'd37: pixel <= 24'h4A_24_FF;
                10'd38: pixel <= 24'h24_FF_EE;
                10'd39: pixel <= 24'hFF_EF_4A;
                10'd40: pixel <= 24'hF1_4B_24;
                10'd41: pixel <= 24'h4B_25_FF;
                10'd42: pixel <= 24'h24_FF_F0;
                10'd43: pixel <= 24'hFF_F1_4B;
                10'd44: pixel <= 24'hF0_4B_25;
                10'd45: pixel <= 24'h4B_24_FF;
                10'd46: pixel <= 24'h25_FF_F0;
                10'd47: pixel <= 24'hFF_F0_4B;
                10'd48: pixel <= 24'hF0_4B_25;
                10'd49: pixel <= 24'h4B_24_FF;
                10'd50: pixel <= 24'h24_FF_EE;
                10'd51: pixel <= 24'hFF_ED_4B;
                10'd52: pixel <= 24'hF2_63_23;
                10'd53: pixel <= 24'h33_3C_FF;
                10'd54: pixel <= 24'h52_FF_A4;
                10'd55: pixel <= 24'hFF_1C_22;
                10'd56: pixel <= 24'h19_19_27;
                10'd57: pixel <= 24'hB2_1F_FF;
                10'd58: pixel <= 24'h1A_FF_FE;
                10'd59: pixel <= 24'hFF_F9_A2;
                10'd60: pixel <= 24'hFB_A1_1C;
                10'd61: pixel <= 24'hA1_1A_FF;
                10'd62: pixel <= 24'h19_FF_FB;
                10'd63: pixel <= 24'hFF_F9_A2;
                10'd64: pixel <= 24'hE8_A9_3F;
                10'd65: pixel <= 24'h22_52_FF;
                10'd66: pixel <= 24'h51_FF_1C;
                10'd67: pixel <= 24'hFF_1C_22;
                10'd68: pixel <= 24'h1D_22_51;
                10'd69: pixel <= 24'h22_51_FF;
                10'd70: pixel <= 24'h51_FF_1D;
                10'd71: pixel <= 24'hFF_1D_23;
                10'd72: pixel <= 24'h52_AF_44;
                10'd73: pixel <= 24'h95_46_FF;
                10'd74: pixel <= 24'h46_FF_18;
                10'd75: pixel <= 24'hFF_18_95;
                10'd76: pixel <= 24'h18_95_47;
                10'd77: pixel <= 24'h95_46_FF;
                10'd78: pixel <= 24'h4C_FF_18;
                10'd79: pixel <= 24'hFF_48_B1;
                10'd80: pixel <= 24'h1D_23_52;
                10'd81: pixel <= 24'h22_51_FF;
                10'd82: pixel <= 24'h52_FF_20;
                10'd83: pixel <= 24'hFF_1D_23;
                10'd84: pixel <= 24'h1D_23_52;
                10'd85: pixel <= 24'h23_52_FF;
                10'd86: pixel <= 24'h53_FF_1D;
                10'd87: pixel <= 24'hFF_1D_23;
                10'd88: pixel <= 24'h11_29_37;
                10'd89: pixel <= 24'hB2_4F_FF;
                10'd90: pixel <= 24'h4D_FF_3A;
                10'd91: pixel <= 24'hFF_19_94;
                10'd92: pixel <= 24'h1F_83_3B;
                10'd93: pixel <= 24'h21_50_FF;
                10'd94: pixel <= 24'hD7_FF_1D;
                10'd95: pixel <= 24'hFF_0A_A2;
                10'd96: pixel <= 24'h20_7F_C2;
                10'd97: pixel <= 24'h7F_C2_FF;
                10'd98: pixel <= 24'hC2_FF_1F;
                10'd99: pixel <= 24'hFF_1F_7F;
            endcase
            10'd17: case (x)
                10'd0: pixel <= 24'h93_77_41;
                10'd1: pixel <= 24'hA1_2E_FF;
                10'd2: pixel <= 24'h20_FF_FC;
                10'd3: pixel <= 24'hFF_EF_6E;
                10'd4: pixel <= 24'hEF_6F_21;
                10'd5: pixel <= 24'h6E_21_FF;
                10'd6: pixel <= 24'h22_FF_F1;
                10'd7: pixel <= 24'hFF_F3_6C;
                10'd8: pixel <= 24'hF1_6D_22;
                10'd9: pixel <= 24'h6E_24_FF;
                10'd10: pixel <= 24'h24_FF_F4;
                10'd11: pixel <= 24'hFF_F3_6E;
                10'd12: pixel <= 24'hF3_6E_24;
                10'd13: pixel <= 24'h6D_24_FF;
                10'd14: pixel <= 24'h25_FF_F3;
                10'd15: pixel <= 24'hFF_F4_6D;
                10'd16: pixel <= 24'hF3_6D_26;
                10'd17: pixel <= 24'h6D_26_FF;
                10'd18: pixel <= 24'h29_FF_F3;
                10'd19: pixel <= 24'hFF_F6_6E;
                10'd20: pixel <= 24'hF6_5F_2F;
                10'd21: pixel <= 24'h24_55_FF;
                10'd22: pixel <= 24'h29_FF_20;
                10'd23: pixel <= 24'hFF_1A_1C;
                10'd24: pixel <= 24'hF6_B5_18;
                10'd25: pixel <= 24'hB4_1A_FF;
                10'd26: pixel <= 24'h18_FF_F7;
                10'd27: pixel <= 24'hFF_F7_B4;
                10'd28: pixel <= 24'hF7_B5_16;
                10'd29: pixel <= 24'hB4_15_FF;
                10'd30: pixel <= 24'h3D_FF_FB;
                10'd31: pixel <= 24'hFF_E5_A7;
                10'd32: pixel <= 24'h20_23_54;
                10'd33: pixel <= 24'h24_54_FF;
                10'd34: pixel <= 24'h54_FF_1E;
                10'd35: pixel <= 24'hFF_20_23;
                10'd36: pixel <= 24'h20_23_54;
                10'd37: pixel <= 24'h24_54_FF;
                10'd38: pixel <= 24'h42_FF_1E;
                10'd39: pixel <= 24'hFF_51_AE;
                10'd40: pixel <= 24'h3F_B0_4B;
                10'd41: pixel <= 24'hB3_47_FF;
                10'd42: pixel <= 24'h49_FF_3E;
                10'd43: pixel <= 24'hFF_3E_B2;
                10'd44: pixel <= 24'h3C_B3_47;
                10'd45: pixel <= 24'hB1_47_FF;
                10'd46: pixel <= 24'h53_FF_4A;
                10'd47: pixel <= 24'hFF_1B_23;
                10'd48: pixel <= 24'h21_22_54;
                10'd49: pixel <= 24'h24_54_FF;
                10'd50: pixel <= 24'h54_FF_1E;
                10'd51: pixel <= 24'hFF_1E_24;
                10'd52: pixel <= 24'h1E_24_54;
                10'd53: pixel <= 24'h24_54_FF;
                10'd54: pixel <= 24'h54_FF_1E;
                10'd55: pixel <= 24'hFF_1F_23;
                10'd56: pixel <= 24'h30_8D_4C;
                10'd57: pixel <= 24'hB5_4B_FF;
                10'd58: pixel <= 24'h37_FF_3A;
                10'd59: pixel <= 24'hFF_1C_82;
                10'd60: pixel <= 24'h1D_23_4F;
                10'd61: pixel <= 24'h9E_CE_FF;
                10'd62: pixel <= 24'hDD_FF_06;
                10'd63: pixel <= 24'hFF_0A_A5;
                10'd64: pixel <= 24'h09_A5_DE;
                10'd65: pixel <= 24'hA4_DF_FF;
                10'd66: pixel <= 24'hDA_FF_0A;
                10'd67: pixel <= 24'hFF_0B_A4;
                10'd68: pixel <= 24'h18_7E_C2;
                10'd69: pixel <= 24'h25_52_FF;
                10'd70: pixel <= 24'hA2_FF_1C;
                10'd71: pixel <= 24'hFF_B7_50;
                10'd72: pixel <= 24'h9F_2B_8A;
                10'd73: pixel <= 24'h2C_8D_FF;
                10'd74: pixel <= 24'h8D_FF_9D;
                10'd75: pixel <= 24'hFF_9C_2C;
                10'd76: pixel <= 24'h9D_2C_8D;
                10'd77: pixel <= 24'h2C_8E_FF;
                10'd78: pixel <= 24'h8E_FF_9D;
                10'd79: pixel <= 24'hFF_9D_2C;
                10'd80: pixel <= 24'h9D_2C_8E;
                10'd81: pixel <= 24'h2C_8E_FF;
                10'd82: pixel <= 24'h8E_FF_9C;
                10'd83: pixel <= 24'hFF_9A_2D;
                10'd84: pixel <= 24'h86_29_7E;
                10'd85: pixel <= 24'h29_69_FF;
                10'd86: pixel <= 24'h51_FF_5B;
                10'd87: pixel <= 24'hFF_1D_23;
                10'd88: pixel <= 24'h1E_22_53;
                10'd89: pixel <= 24'h22_53_FF;
                10'd90: pixel <= 24'h53_FF_1E;
                10'd91: pixel <= 24'hFF_1D_23;
                10'd92: pixel <= 24'h1D_23_53;
                10'd93: pixel <= 24'h25_50_FF;
                10'd94: pixel <= 24'h9E_FF_1C;
                10'd95: pixel <= 24'hFF_33_58;
                10'd96: pixel <= 24'h30_59_A0;
                10'd97: pixel <= 24'h5A_9F_FF;
                10'd98: pixel <= 24'h81_FF_30;
                10'd99: pixel <= 24'hFF_22_41;
            endcase
            10'd18: case (x)
                10'd0: pixel <= 24'h21_24_55;
                10'd1: pixel <= 24'h24_55_FF;
                10'd2: pixel <= 24'h55_FF_21;
                10'd3: pixel <= 24'hFF_21_24;
                10'd4: pixel <= 24'h20_24_57;
                10'd5: pixel <= 24'h24_55_FF;
                10'd6: pixel <= 24'h56_FF_21;
                10'd7: pixel <= 24'hFF_20_24;
                10'd8: pixel <= 24'h21_23_58;
                10'd9: pixel <= 24'h23_58_FF;
                10'd10: pixel <= 24'h56_FF_22;
                10'd11: pixel <= 24'hFF_20_24;
                10'd12: pixel <= 24'h21_24_58;
                10'd13: pixel <= 24'h25_56_FF;
                10'd14: pixel <= 24'h55_FF_20;
                10'd15: pixel <= 24'hFF_22_23;
                10'd16: pixel <= 24'h1F_25_55;
                10'd17: pixel <= 24'h24_55_FF;
                10'd18: pixel <= 24'h55_FF_21;
                10'd19: pixel <= 24'hFF_21_24;
                10'd20: pixel <= 24'h1F_25_55;
                10'd21: pixel <= 24'h25_55_FF;
                10'd22: pixel <= 24'h56_FF_1F;
                10'd23: pixel <= 24'hFF_20_24;
                10'd24: pixel <= 24'h21_23_5A;
                10'd25: pixel <= 24'h25_57_FF;
                10'd26: pixel <= 24'h53_FF_20;
                10'd27: pixel <= 24'hFF_20_23;
                10'd28: pixel <= 24'h1F_24_5A;
                10'd29: pixel <= 24'h24_58_FF;
                10'd30: pixel <= 24'h58_FF_20;
                10'd31: pixel <= 24'hFF_1E_25;
                10'd32: pixel <= 24'h20_25_56;
                10'd33: pixel <= 24'h25_52_FF;
                10'd34: pixel <= 24'h57_FF_21;
                10'd35: pixel <= 24'hFF_23_23;
                10'd36: pixel <= 24'h21_24_56;
                10'd37: pixel <= 24'h23_56_FF;
                10'd38: pixel <= 24'h53_FF_22;
                10'd39: pixel <= 24'hFF_21_25;
                10'd40: pixel <= 24'h21_24_55;
                10'd41: pixel <= 24'h25_57_FF;
                10'd42: pixel <= 24'h55_FF_20;
                10'd43: pixel <= 24'hFF_1E_26;
                10'd44: pixel <= 24'h1E_25_56;
                10'd45: pixel <= 24'h25_56_FF;
                10'd46: pixel <= 24'h57_FF_20;
                10'd47: pixel <= 24'hFF_20_25;
                10'd48: pixel <= 24'h20_25_56;
                10'd49: pixel <= 24'h25_56_FF;
                10'd50: pixel <= 24'h56_FF_1F;
                10'd51: pixel <= 24'hFF_20_25;
                10'd52: pixel <= 24'h21_24_55;
                10'd53: pixel <= 24'h24_55_FF;
                10'd54: pixel <= 24'h55_FF_21;
                10'd55: pixel <= 24'hFF_1F_25;
                10'd56: pixel <= 24'h1F_25_55;
                10'd57: pixel <= 24'h24_55_FF;
                10'd58: pixel <= 24'h55_FF_21;
                10'd59: pixel <= 24'hFF_21_24;
                10'd60: pixel <= 24'h1C_25_50;
                10'd61: pixel <= 24'h58_9F_FF;
                10'd62: pixel <= 24'hA1_FF_36;
                10'd63: pixel <= 24'hFF_31_5A;
                10'd64: pixel <= 24'h31_5A_A1;
                10'd65: pixel <= 24'h41_81_FF;
                10'd66: pixel <= 24'h81_FF_22;
                10'd67: pixel <= 24'hFF_22_41;
                10'd68: pixel <= 24'h30_59_A0;
                10'd69: pixel <= 24'h59_A0_FF;
                10'd70: pixel <= 24'h9F_FF_30;
                10'd71: pixel <= 24'hFF_35_59;
                10'd72: pixel <= 24'h1A_2A_5E;
                10'd73: pixel <= 24'h24_52_FF;
                10'd74: pixel <= 24'h54_FF_1E;
                10'd75: pixel <= 24'hFF_1E_24;
                10'd76: pixel <= 24'h1E_24_54;
                10'd77: pixel <= 24'h23_54_FF;
                10'd78: pixel <= 24'h54_FF_20;
                10'd79: pixel <= 24'hFF_1E_24;
                10'd80: pixel <= 24'h1E_24_54;
                10'd81: pixel <= 24'h1F_4C_FF;
                10'd82: pixel <= 24'h36_FF_20;
                10'd83: pixel <= 24'hFF_EC_24;
                10'd84: pixel <= 24'hEF_23_34;
                10'd85: pixel <= 24'h23_35_FF;
                10'd86: pixel <= 24'h38_FF_EF;
                10'd87: pixel <= 24'hFF_EC_23;
                10'd88: pixel <= 24'hEE_23_36;
                10'd89: pixel <= 24'h29_38_FF;
                10'd90: pixel <= 24'h54_FF_ED;
                10'd91: pixel <= 24'hFF_20_23;
                10'd92: pixel <= 24'h1E_24_54;
                10'd93: pixel <= 24'h24_54_FF;
                10'd94: pixel <= 24'h54_FF_1E;
                10'd95: pixel <= 24'hFF_1E_24;
                10'd96: pixel <= 24'h20_23_54;
                10'd97: pixel <= 24'h23_54_FF;
                10'd98: pixel <= 24'h54_FF_20;
                10'd99: pixel <= 24'hFF_21_24;
            endcase
            10'd19: case (x)
                10'd0: pixel <= 24'h22_25_58;
                10'd1: pixel <= 24'h25_58_FF;
                10'd2: pixel <= 24'h58_FF_22;
                10'd3: pixel <= 24'hFF_22_25;
                10'd4: pixel <= 24'h22_25_58;
                10'd5: pixel <= 24'h25_58_FF;
                10'd6: pixel <= 24'h58_FF_22;
                10'd7: pixel <= 24'hFF_20_26;
                10'd8: pixel <= 24'h22_25_58;
                10'd9: pixel <= 24'h25_58_FF;
                10'd10: pixel <= 24'h58_FF_22;
                10'd11: pixel <= 24'hFF_22_25;
                10'd12: pixel <= 24'h22_25_58;
                10'd13: pixel <= 24'h25_58_FF;
                10'd14: pixel <= 24'h58_FF_22;
                10'd15: pixel <= 24'hFF_22_25;
                10'd16: pixel <= 24'h22_25_58;
                10'd17: pixel <= 24'h25_58_FF;
                10'd18: pixel <= 24'h58_FF_22;
                10'd19: pixel <= 24'hFF_22_25;
                10'd20: pixel <= 24'h22_25_58;
                10'd21: pixel <= 24'h25_58_FF;
                10'd22: pixel <= 24'h58_FF_22;
                10'd23: pixel <= 24'hFF_22_25;
                10'd24: pixel <= 24'h22_25_58;
                10'd25: pixel <= 24'h26_58_FF;
                10'd26: pixel <= 24'h51_FF_20;
                10'd27: pixel <= 24'hFF_1E_27;
                10'd28: pixel <= 24'h35_59_9F;
                10'd29: pixel <= 24'h5B_A4_FF;
                10'd30: pixel <= 24'hA3_FF_33;
                10'd31: pixel <= 24'hFF_34_5D;
                10'd32: pixel <= 24'h22_41_81;
                10'd33: pixel <= 24'h40_81_FF;
                10'd34: pixel <= 24'hA1_FF_24;
                10'd35: pixel <= 24'hFF_31_5A;
                10'd36: pixel <= 24'h31_5A_A1;
                10'd37: pixel <= 24'h5A_A0_FF;
                10'd38: pixel <= 24'h5E_FF_36;
                10'd39: pixel <= 24'hFF_18_2B;
                10'd40: pixel <= 24'h21_24_55;
                10'd41: pixel <= 24'h25_55_FF;
                10'd42: pixel <= 24'h55_FF_1F;
                10'd43: pixel <= 24'hFF_21_24;
                10'd44: pixel <= 24'h1F_25_55;
                10'd45: pixel <= 24'h24_55_FF;
                10'd46: pixel <= 24'h55_FF_21;
                10'd47: pixel <= 24'hFF_1F_25;
                10'd48: pixel <= 24'h1F_25_56;
                10'd49: pixel <= 24'h25_54_FF;
                10'd50: pixel <= 24'h56_FF_1F;
                10'd51: pixel <= 24'hFF_22_23;
                10'd52: pixel <= 24'h20_24_55;
                10'd53: pixel <= 24'h24_56_FF;
                10'd54: pixel <= 24'h56_FF_20;
                10'd55: pixel <= 24'hFF_25_22;
                10'd56: pixel <= 24'h22_23_57;
                10'd57: pixel <= 24'h24_55_FF;
                10'd58: pixel <= 24'h55_FF_21;
                10'd59: pixel <= 24'hFF_21_24;
                10'd60: pixel <= 24'h21_24_55;
                10'd61: pixel <= 24'h25_55_FF;
                10'd62: pixel <= 24'h55_FF_1F;
                10'd63: pixel <= 24'hFF_1F_25;
                10'd64: pixel <= 24'h1F_25_55;
                10'd65: pixel <= 24'h25_55_FF;
                10'd66: pixel <= 24'h57_FF_1F;
                10'd67: pixel <= 24'hFF_1F_25;
                10'd68: pixel <= 24'h1F_23_53;
                10'd69: pixel <= 24'h26_56_FF;
                10'd70: pixel <= 24'h56_FF_1F;
                10'd71: pixel <= 24'hFF_24_24;
                10'd72: pixel <= 24'h20_24_56;
                10'd73: pixel <= 24'h23_58_FF;
                10'd74: pixel <= 24'h58_FF_21;
                10'd75: pixel <= 24'hFF_20_24;
                10'd76: pixel <= 24'h1D_24_55;
                10'd77: pixel <= 24'h23_56_FF;
                10'd78: pixel <= 24'h57_FF_20;
                10'd79: pixel <= 24'hFF_20_22;
                10'd80: pixel <= 24'h1E_23_56;
                10'd81: pixel <= 24'h24_55_FF;
                10'd82: pixel <= 24'h55_FF_1D;
                10'd83: pixel <= 24'hFF_1E_23;
                10'd84: pixel <= 24'h20_22_57;
                10'd85: pixel <= 24'h22_57_FF;
                10'd86: pixel <= 24'h56_FF_21;
                10'd87: pixel <= 24'hFF_1F_23;
                10'd88: pixel <= 24'h1F_23_55;
                10'd89: pixel <= 24'h23_53_FF;
                10'd90: pixel <= 24'h54_FF_21;
                10'd91: pixel <= 24'hFF_20_23;
                10'd92: pixel <= 24'h20_23_56;
                10'd93: pixel <= 24'h23_56_FF;
                10'd94: pixel <= 24'h58_FF_20;
                10'd95: pixel <= 24'hFF_20_22;
                10'd96: pixel <= 24'h1F_23_58;
                10'd97: pixel <= 24'h22_51_FF;
                10'd98: pixel <= 24'h54_FF_23;
                10'd99: pixel <= 24'hFF_20_23;
            endcase
            10'd20: case (x)
                10'd0: pixel <= 24'h22_41_81;
                10'd1: pixel <= 24'h5B_A4_FF;
                10'd2: pixel <= 24'hA4_FF_33;
                10'd3: pixel <= 24'hFF_33_5B;
                10'd4: pixel <= 24'h37_5B_A3;
                10'd5: pixel <= 24'h2C_61_FF;
                10'd6: pixel <= 24'h58_FF_19;
                10'd7: pixel <= 24'hFF_20_26;
                10'd8: pixel <= 24'h22_25_58;
                10'd9: pixel <= 24'h25_58_FF;
                10'd10: pixel <= 24'h58_FF_22;
                10'd11: pixel <= 24'hFF_22_25;
                10'd12: pixel <= 24'h20_26_58;
                10'd13: pixel <= 24'h25_58_FF;
                10'd14: pixel <= 24'h58_FF_22;
                10'd15: pixel <= 24'hFF_22_25;
                10'd16: pixel <= 24'h22_25_58;
                10'd17: pixel <= 24'h25_58_FF;
                10'd18: pixel <= 24'h58_FF_22;
                10'd19: pixel <= 24'hFF_20_26;
                10'd20: pixel <= 24'h22_25_58;
                10'd21: pixel <= 24'h26_58_FF;
                10'd22: pixel <= 24'h58_FF_20;
                10'd23: pixel <= 24'hFF_22_25;
                10'd24: pixel <= 24'h20_26_58;
                10'd25: pixel <= 24'h25_58_FF;
                10'd26: pixel <= 24'h58_FF_22;
                10'd27: pixel <= 24'hFF_22_25;
                10'd28: pixel <= 24'h22_25_58;
                10'd29: pixel <= 24'h25_58_FF;
                10'd30: pixel <= 24'h58_FF_22;
                10'd31: pixel <= 24'hFF_22_25;
                10'd32: pixel <= 24'h22_25_58;
                10'd33: pixel <= 24'h25_58_FF;
                10'd34: pixel <= 24'h58_FF_22;
                10'd35: pixel <= 24'hFF_22_25;
                10'd36: pixel <= 24'h22_25_58;
                10'd37: pixel <= 24'h25_58_FF;
                10'd38: pixel <= 24'h58_FF_22;
                10'd39: pixel <= 24'hFF_22_25;
                10'd40: pixel <= 24'h20_26_58;
                10'd41: pixel <= 24'h25_58_FF;
                10'd42: pixel <= 24'h58_FF_22;
                10'd43: pixel <= 24'hFF_22_25;
                10'd44: pixel <= 24'h22_25_58;
                10'd45: pixel <= 24'h25_58_FF;
                10'd46: pixel <= 24'h58_FF_22;
                10'd47: pixel <= 24'hFF_22_25;
                10'd48: pixel <= 24'h22_25_58;
                10'd49: pixel <= 24'h25_58_FF;
                10'd50: pixel <= 24'h58_FF_22;
                10'd51: pixel <= 24'hFF_22_25;
                10'd52: pixel <= 24'h20_26_58;
                10'd53: pixel <= 24'h25_58_FF;
                10'd54: pixel <= 24'h58_FF_22;
                10'd55: pixel <= 24'hFF_22_25;
                10'd56: pixel <= 24'h22_25_58;
                10'd57: pixel <= 24'h26_58_FF;
                10'd58: pixel <= 24'h58_FF_20;
                10'd59: pixel <= 24'hFF_20_26;
                10'd60: pixel <= 24'h22_25_58;
                10'd61: pixel <= 24'h25_58_FF;
                10'd62: pixel <= 24'h58_FF_22;
                10'd63: pixel <= 24'hFF_22_25;
                10'd64: pixel <= 24'h22_25_58;
                10'd65: pixel <= 24'h25_58_FF;
                10'd66: pixel <= 24'h58_FF_22;
                10'd67: pixel <= 24'hFF_20_26;
                10'd68: pixel <= 24'h22_25_58;
                10'd69: pixel <= 24'h25_58_FF;
                10'd70: pixel <= 24'h58_FF_22;
                10'd71: pixel <= 24'hFF_20_26;
                10'd72: pixel <= 24'h22_25_58;
                10'd73: pixel <= 24'h26_58_FF;
                10'd74: pixel <= 24'h58_FF_20;
                10'd75: pixel <= 24'hFF_22_25;
                10'd76: pixel <= 24'h20_26_58;
                10'd77: pixel <= 24'h25_58_FF;
                10'd78: pixel <= 24'h58_FF_22;
                10'd79: pixel <= 24'hFF_22_25;
                10'd80: pixel <= 24'h22_25_58;
                10'd81: pixel <= 24'h25_58_FF;
                10'd82: pixel <= 24'h58_FF_22;
                10'd83: pixel <= 24'hFF_22_25;
                10'd84: pixel <= 24'h22_25_58;
                10'd85: pixel <= 24'h26_58_FF;
                10'd86: pixel <= 24'h58_FF_20;
                10'd87: pixel <= 24'hFF_22_25;
                10'd88: pixel <= 24'h22_25_58;
                10'd89: pixel <= 24'h25_58_FF;
                10'd90: pixel <= 24'h58_FF_22;
                10'd91: pixel <= 24'hFF_22_25;
                10'd92: pixel <= 24'h22_25_58;
                10'd93: pixel <= 24'h25_58_FF;
                10'd94: pixel <= 24'h58_FF_22;
                10'd95: pixel <= 24'hFF_22_25;
                10'd96: pixel <= 24'h22_25_58;
                10'd97: pixel <= 24'h25_58_FF;
                10'd98: pixel <= 24'h58_FF_22;
                10'd99: pixel <= 24'hFF_22_25;
            endcase
            10'd21: case (x)
                10'd0: pixel <= 24'h20_26_58;
                10'd1: pixel <= 24'h25_58_FF;
                10'd2: pixel <= 24'h58_FF_22;
                10'd3: pixel <= 24'hFF_20_26;
                10'd4: pixel <= 24'h20_26_58;
                10'd5: pixel <= 24'h25_5A_FF;
                10'd6: pixel <= 24'h58_FF_22;
                10'd7: pixel <= 24'hFF_20_26;
                10'd8: pixel <= 24'h22_25_58;
                10'd9: pixel <= 24'h26_58_FF;
                10'd10: pixel <= 24'h5A_FF_20;
                10'd11: pixel <= 24'hFF_22_25;
                10'd12: pixel <= 24'h20_26_58;
                10'd13: pixel <= 24'h26_58_FF;
                10'd14: pixel <= 24'h58_FF_20;
                10'd15: pixel <= 24'hFF_20_26;
                10'd16: pixel <= 24'h20_26_58;
                10'd17: pixel <= 24'h25_5A_FF;
                10'd18: pixel <= 24'h58_FF_20;
                10'd19: pixel <= 24'hFF_20_26;
                10'd20: pixel <= 24'h20_26_58;
                10'd21: pixel <= 24'h26_58_FF;
                10'd22: pixel <= 24'h5A_FF_20;
                10'd23: pixel <= 24'hFF_20_25;
                10'd24: pixel <= 24'h20_26_58;
                10'd25: pixel <= 24'h26_58_FF;
                10'd26: pixel <= 24'h58_FF_20;
                10'd27: pixel <= 24'hFF_20_26;
                10'd28: pixel <= 24'h20_26_58;
                10'd29: pixel <= 24'h26_58_FF;
                10'd30: pixel <= 24'h58_FF_20;
                10'd31: pixel <= 24'hFF_20_26;
                10'd32: pixel <= 24'h20_25_5A;
                10'd33: pixel <= 24'h26_58_FF;
                10'd34: pixel <= 24'h58_FF_20;
                10'd35: pixel <= 24'hFF_20_26;
                10'd36: pixel <= 24'h20_26_58;
                10'd37: pixel <= 24'h26_58_FF;
                10'd38: pixel <= 24'h58_FF_20;
                10'd39: pixel <= 24'hFF_20_26;
                10'd40: pixel <= 24'h20_26_58;
                10'd41: pixel <= 24'h26_58_FF;
                10'd42: pixel <= 24'h58_FF_20;
                10'd43: pixel <= 24'hFF_20_26;
                10'd44: pixel <= 24'h20_26_58;
                10'd45: pixel <= 24'h26_58_FF;
                10'd46: pixel <= 24'h58_FF_20;
                10'd47: pixel <= 24'hFF_20_26;
                10'd48: pixel <= 24'h20_26_58;
                10'd49: pixel <= 24'h26_58_FF;
                10'd50: pixel <= 24'h58_FF_20;
                10'd51: pixel <= 24'hFF_20_26;
                10'd52: pixel <= 24'h20_26_58;
                10'd53: pixel <= 24'h26_58_FF;
                10'd54: pixel <= 24'h58_FF_20;
                10'd55: pixel <= 24'hFF_20_26;
                10'd56: pixel <= 24'h20_26_58;
                10'd57: pixel <= 24'h26_58_FF;
                10'd58: pixel <= 24'h58_FF_20;
                10'd59: pixel <= 24'hFF_20_26;
                10'd60: pixel <= 24'h20_26_58;
                10'd61: pixel <= 24'h26_58_FF;
                10'd62: pixel <= 24'h58_FF_20;
                10'd63: pixel <= 24'hFF_20_26;
                10'd64: pixel <= 24'h20_26_58;
                10'd65: pixel <= 24'h26_58_FF;
                10'd66: pixel <= 24'h58_FF_20;
                10'd67: pixel <= 24'hFF_20_26;
                10'd68: pixel <= 24'h20_26_58;
                10'd69: pixel <= 24'h26_58_FF;
                10'd70: pixel <= 24'h58_FF_20;
                10'd71: pixel <= 24'hFF_20_26;
                10'd72: pixel <= 24'h20_26_58;
                10'd73: pixel <= 24'h26_58_FF;
                10'd74: pixel <= 24'h58_FF_20;
                10'd75: pixel <= 24'hFF_20_26;
                10'd76: pixel <= 24'h20_26_58;
                10'd77: pixel <= 24'h26_58_FF;
                10'd78: pixel <= 24'h58_FF_20;
                10'd79: pixel <= 24'hFF_20_26;
                10'd80: pixel <= 24'h20_26_58;
                10'd81: pixel <= 24'h26_58_FF;
                10'd82: pixel <= 24'h58_FF_20;
                10'd83: pixel <= 24'hFF_20_26;
                10'd84: pixel <= 24'h20_25_5A;
                10'd85: pixel <= 24'h26_58_FF;
                10'd86: pixel <= 24'h58_FF_20;
                10'd87: pixel <= 24'hFF_20_26;
                10'd88: pixel <= 24'h20_26_58;
                10'd89: pixel <= 24'h26_58_FF;
                10'd90: pixel <= 24'h58_FF_20;
                10'd91: pixel <= 24'hFF_20_26;
                10'd92: pixel <= 24'h20_26_58;
                10'd93: pixel <= 24'h26_55_FF;
                10'd94: pixel <= 24'hA2_FF_1E;
                10'd95: pixel <= 24'hFF_38_5D;
                10'd96: pixel <= 24'h34_5C_A5;
                10'd97: pixel <= 24'h5D_A3_FF;
                10'd98: pixel <= 24'h81_FF_34;
                10'd99: pixel <= 24'hFF_22_41;
            endcase
            10'd22: case (x)
                10'd0: pixel <= 24'h22_27_5B;
                10'd1: pixel <= 24'h27_5B_FF;
                10'd2: pixel <= 24'h5B_FF_22;
                10'd3: pixel <= 24'hFF_22_27;
                10'd4: pixel <= 24'h22_27_5B;
                10'd5: pixel <= 24'h27_5B_FF;
                10'd6: pixel <= 24'h5B_FF_22;
                10'd7: pixel <= 24'hFF_22_27;
                10'd8: pixel <= 24'h22_27_5B;
                10'd9: pixel <= 24'h27_5B_FF;
                10'd10: pixel <= 24'h5B_FF_22;
                10'd11: pixel <= 24'hFF_22_27;
                10'd12: pixel <= 24'h22_27_5B;
                10'd13: pixel <= 24'h27_5B_FF;
                10'd14: pixel <= 24'h5B_FF_22;
                10'd15: pixel <= 24'hFF_22_27;
                10'd16: pixel <= 24'h22_27_5B;
                10'd17: pixel <= 24'h27_5B_FF;
                10'd18: pixel <= 24'h5B_FF_22;
                10'd19: pixel <= 24'hFF_22_27;
                10'd20: pixel <= 24'h29_37_74;
                10'd21: pixel <= 24'h39_75_FF;
                10'd22: pixel <= 24'h72_FF_25;
                10'd23: pixel <= 24'hFF_24_37;
                10'd24: pixel <= 24'h24_36_72;
                10'd25: pixel <= 24'h36_72_FF;
                10'd26: pixel <= 24'h71_FF_24;
                10'd27: pixel <= 24'hFF_23_35;
                10'd28: pixel <= 24'h21_32_6F;
                10'd29: pixel <= 24'h33_6D_FF;
                10'd30: pixel <= 24'h6B_FF_21;
                10'd31: pixel <= 24'hFF_20_32;
                10'd32: pixel <= 24'h20_32_6B;
                10'd33: pixel <= 24'h2F_67_FF;
                10'd34: pixel <= 24'h67_FF_1D;
                10'd35: pixel <= 24'hFF_1C_2E;
                10'd36: pixel <= 24'h1C_2E_67;
                10'd37: pixel <= 24'h2C_66_FF;
                10'd38: pixel <= 24'h63_FF_1D;
                10'd39: pixel <= 24'hFF_1B_2E;
                10'd40: pixel <= 24'h1A_2B_5F;
                10'd41: pixel <= 24'h2C_5F_FF;
                10'd42: pixel <= 24'h5B_FF_19;
                10'd43: pixel <= 24'hFF_18_29;
                10'd44: pixel <= 24'h17_28_5A;
                10'd45: pixel <= 24'h28_58_FF;
                10'd46: pixel <= 24'h54_FF_17;
                10'd47: pixel <= 24'hFF_17_27;
                10'd48: pixel <= 24'h17_28_52;
                10'd49: pixel <= 24'h24_52_FF;
                10'd50: pixel <= 24'h50_FF_16;
                10'd51: pixel <= 24'hFF_15_24;
                10'd52: pixel <= 24'h15_23_4F;
                10'd53: pixel <= 24'h21_4D_FF;
                10'd54: pixel <= 24'h4E_FF_14;
                10'd55: pixel <= 24'hFF_14_22;
                10'd56: pixel <= 24'h12_1F_4B;
                10'd57: pixel <= 24'h1F_4B_FF;
                10'd58: pixel <= 24'h4A_FF_12;
                10'd59: pixel <= 24'hFF_12_1D;
                10'd60: pixel <= 24'h10_1E_47;
                10'd61: pixel <= 24'h60_A8_FF;
                10'd62: pixel <= 24'hA9_FF_3B;
                10'd63: pixel <= 24'hFF_37_60;
                10'd64: pixel <= 24'h36_5F_A5;
                10'd65: pixel <= 24'h41_81_FF;
                10'd66: pixel <= 24'h81_FF_22;
                10'd67: pixel <= 24'hFF_24_40;
                10'd68: pixel <= 24'h34_5C_A5;
                10'd69: pixel <= 24'h5D_A6_FF;
                10'd70: pixel <= 24'hA5_FF_35;
                10'd71: pixel <= 24'hFF_39_5D;
                10'd72: pixel <= 24'h1A_2D_62;
                10'd73: pixel <= 24'h26_58_FF;
                10'd74: pixel <= 24'h5A_FF_20;
                10'd75: pixel <= 24'hFF_20_25;
                10'd76: pixel <= 24'h20_26_58;
                10'd77: pixel <= 24'h26_58_FF;
                10'd78: pixel <= 24'h58_FF_20;
                10'd79: pixel <= 24'hFF_20_26;
                10'd80: pixel <= 24'h20_25_5A;
                10'd81: pixel <= 24'h26_58_FF;
                10'd82: pixel <= 24'h58_FF_20;
                10'd83: pixel <= 24'hFF_20_26;
                10'd84: pixel <= 24'h20_25_5A;
                10'd85: pixel <= 24'h26_58_FF;
                10'd86: pixel <= 24'h58_FF_20;
                10'd87: pixel <= 24'hFF_20_26;
                10'd88: pixel <= 24'h20_26_58;
                10'd89: pixel <= 24'h26_58_FF;
                10'd90: pixel <= 24'h58_FF_20;
                10'd91: pixel <= 24'hFF_20_26;
                10'd92: pixel <= 24'h20_26_58;
                10'd93: pixel <= 24'h26_58_FF;
                10'd94: pixel <= 24'h58_FF_20;
                10'd95: pixel <= 24'hFF_20_26;
                10'd96: pixel <= 24'h22_25_58;
                10'd97: pixel <= 24'h26_58_FF;
                10'd98: pixel <= 24'h58_FF_20;
                10'd99: pixel <= 24'hFF_20_26;
            endcase
            10'd23: case (x)
                10'd0: pixel <= 24'h37_60_A9;
                10'd1: pixel <= 24'h60_A9_FF;
                10'd2: pixel <= 24'hA9_FF_37;
                10'd3: pixel <= 24'hFF_37_60;
                10'd4: pixel <= 24'h37_60_A9;
                10'd5: pixel <= 24'h60_A9_FF;
                10'd6: pixel <= 24'hA9_FF_37;
                10'd7: pixel <= 24'hFF_37_60;
                10'd8: pixel <= 24'h37_60_A9;
                10'd9: pixel <= 24'h60_A9_FF;
                10'd10: pixel <= 24'hA9_FF_37;
                10'd11: pixel <= 24'hFF_37_60;
                10'd12: pixel <= 24'h37_60_A9;
                10'd13: pixel <= 24'h60_A9_FF;
                10'd14: pixel <= 24'hA9_FF_37;
                10'd15: pixel <= 24'hFF_37_60;
                10'd16: pixel <= 24'h37_60_A9;
                10'd17: pixel <= 24'h60_A9_FF;
                10'd18: pixel <= 24'hA9_FF_37;
                10'd19: pixel <= 24'hFF_37_60;
                10'd20: pixel <= 24'h37_60_A9;
                10'd21: pixel <= 24'h60_A9_FF;
                10'd22: pixel <= 24'hA9_FF_37;
                10'd23: pixel <= 24'hFF_37_60;
                10'd24: pixel <= 24'h37_60_A9;
                10'd25: pixel <= 24'h60_A9_FF;
                10'd26: pixel <= 24'hA9_FF_37;
                10'd27: pixel <= 24'hFF_37_60;
                10'd28: pixel <= 24'h38_60_A7;
                10'd29: pixel <= 24'h61_AA_FF;
                10'd30: pixel <= 24'hA7_FF_38;
                10'd31: pixel <= 24'hFF_37_60;
                10'd32: pixel <= 24'h22_41_81;
                10'd33: pixel <= 24'h41_81_FF;
                10'd34: pixel <= 24'hA7_FF_22;
                10'd35: pixel <= 24'hFF_36_5F;
                10'd36: pixel <= 24'h36_5F_A7;
                10'd37: pixel <= 24'h5F_A6_FF;
                10'd38: pixel <= 24'hB8_FF_39;
                10'd39: pixel <= 24'hFF_5A_77;
                10'd40: pixel <= 24'h5B_78_B8;
                10'd41: pixel <= 24'h76_B7_FF;
                10'd42: pixel <= 24'hB5_FF_59;
                10'd43: pixel <= 24'hFF_58_75;
                10'd44: pixel <= 24'h57_75_B4;
                10'd45: pixel <= 24'h74_B3_FF;
                10'd46: pixel <= 24'hB3_FF_55;
                10'd47: pixel <= 24'hFF_54_75;
                10'd48: pixel <= 24'h54_73_B2;
                10'd49: pixel <= 24'h71_B1_FF;
                10'd50: pixel <= 24'hB0_FF_54;
                10'd51: pixel <= 24'hFF_53_70;
                10'd52: pixel <= 24'h51_6E_B0;
                10'd53: pixel <= 24'h6E_B0_FF;
                10'd54: pixel <= 24'hB0_FF_51;
                10'd55: pixel <= 24'hFF_4E_6B;
                10'd56: pixel <= 24'h4C_6D_AE;
                10'd57: pixel <= 24'h6A_AF_FF;
                10'd58: pixel <= 24'hAD_FF_4C;
                10'd59: pixel <= 24'hFF_4D_6A;
                10'd60: pixel <= 24'h4C_69_AB;
                10'd61: pixel <= 24'h67_AC_FF;
                10'd62: pixel <= 24'hAC_FF_4A;
                10'd63: pixel <= 24'hFF_4A_67;
                10'd64: pixel <= 24'h49_66_AB;
                10'd65: pixel <= 24'h66_AB_FF;
                10'd66: pixel <= 24'hA8_FF_49;
                10'd67: pixel <= 24'hFF_47_64;
                10'd68: pixel <= 24'h47_64_A8;
                10'd69: pixel <= 24'h64_A8_FF;
                10'd70: pixel <= 24'hA6_FF_47;
                10'd71: pixel <= 24'hFF_45_62;
                10'd72: pixel <= 24'h44_61_A5;
                10'd73: pixel <= 24'h5F_A4_FF;
                10'd74: pixel <= 24'hA6_FF_42;
                10'd75: pixel <= 24'hFF_42_5E;
                10'd76: pixel <= 24'h40_5C_A3;
                10'd77: pixel <= 24'h5C_A3_FF;
                10'd78: pixel <= 24'hA3_FF_40;
                10'd79: pixel <= 24'hFF_3F_5D;
                10'd80: pixel <= 24'h21_27_5A;
                10'd81: pixel <= 24'h27_59_FF;
                10'd82: pixel <= 24'h5B_FF_22;
                10'd83: pixel <= 24'hFF_22_27;
                10'd84: pixel <= 24'h22_27_5B;
                10'd85: pixel <= 24'h27_5B_FF;
                10'd86: pixel <= 24'h5B_FF_22;
                10'd87: pixel <= 24'hFF_22_27;
                10'd88: pixel <= 24'h22_27_5B;
                10'd89: pixel <= 24'h27_5B_FF;
                10'd90: pixel <= 24'h5B_FF_22;
                10'd91: pixel <= 24'hFF_22_27;
                10'd92: pixel <= 24'h22_27_5B;
                10'd93: pixel <= 24'h27_5B_FF;
                10'd94: pixel <= 24'h5B_FF_22;
                10'd95: pixel <= 24'hFF_22_27;
                10'd96: pixel <= 24'h22_27_5B;
                10'd97: pixel <= 24'h27_5B_FF;
                10'd98: pixel <= 24'h5B_FF_22;
                10'd99: pixel <= 24'hFF_22_27;
            endcase
            10'd24: case (x)
                10'd0: pixel <= 24'h24_40_81;
                10'd1: pixel <= 24'h60_A9_FF;
                10'd2: pixel <= 24'hA9_FF_37;
                10'd3: pixel <= 24'hFF_37_60;
                10'd4: pixel <= 24'h38_61_AA;
                10'd5: pixel <= 24'h60_A8_FF;
                10'd6: pixel <= 24'hA9_FF_38;
                10'd7: pixel <= 24'hFF_37_60;
                10'd8: pixel <= 24'h37_60_AA;
                10'd9: pixel <= 24'h60_A9_FF;
                10'd10: pixel <= 24'hA9_FF_37;
                10'd11: pixel <= 24'hFF_37_60;
                10'd12: pixel <= 24'h37_60_A9;
                10'd13: pixel <= 24'h60_AA_FF;
                10'd14: pixel <= 24'hA9_FF_37;
                10'd15: pixel <= 24'hFF_37_60;
                10'd16: pixel <= 24'h37_60_A9;
                10'd17: pixel <= 24'h60_AA_FF;
                10'd18: pixel <= 24'hA9_FF_37;
                10'd19: pixel <= 24'hFF_37_60;
                10'd20: pixel <= 24'h37_60_A9;
                10'd21: pixel <= 24'h60_A9_FF;
                10'd22: pixel <= 24'hA9_FF_37;
                10'd23: pixel <= 24'hFF_37_60;
                10'd24: pixel <= 24'h37_60_A9;
                10'd25: pixel <= 24'h60_A9_FF;
                10'd26: pixel <= 24'hA9_FF_37;
                10'd27: pixel <= 24'hFF_37_60;
                10'd28: pixel <= 24'h37_60_A9;
                10'd29: pixel <= 24'h60_A9_FF;
                10'd30: pixel <= 24'hA9_FF_37;
                10'd31: pixel <= 24'hFF_37_60;
                10'd32: pixel <= 24'h37_60_A9;
                10'd33: pixel <= 24'h60_A9_FF;
                10'd34: pixel <= 24'hA9_FF_37;
                10'd35: pixel <= 24'hFF_37_60;
                10'd36: pixel <= 24'h37_60_A9;
                10'd37: pixel <= 24'h60_A9_FF;
                10'd38: pixel <= 24'hA9_FF_37;
                10'd39: pixel <= 24'hFF_37_60;
                10'd40: pixel <= 24'h37_60_A9;
                10'd41: pixel <= 24'h60_A9_FF;
                10'd42: pixel <= 24'hA9_FF_37;
                10'd43: pixel <= 24'hFF_37_60;
                10'd44: pixel <= 24'h37_60_A8;
                10'd45: pixel <= 24'h42_81_FF;
                10'd46: pixel <= 24'h5D_FF_1F;
                10'd47: pixel <= 24'hFF_24_27;
                10'd48: pixel <= 24'h23_28_5D;
                10'd49: pixel <= 24'h27_5F_FF;
                10'd50: pixel <= 24'h5D_FF_23;
                10'd51: pixel <= 24'hFF_23_28;
                10'd52: pixel <= 24'h23_27_5F;
                10'd53: pixel <= 24'h28_5D_FF;
                10'd54: pixel <= 24'h5F_FF_23;
                10'd55: pixel <= 24'hFF_23_27;
                10'd56: pixel <= 24'h23_28_5D;
                10'd57: pixel <= 24'h27_5F_FF;
                10'd58: pixel <= 24'h5F_FF_23;
                10'd59: pixel <= 24'hFF_23_27;
                10'd60: pixel <= 24'h23_28_5D;
                10'd61: pixel <= 24'h27_5F_FF;
                10'd62: pixel <= 24'h5D_FF_23;
                10'd63: pixel <= 24'hFF_23_28;
                10'd64: pixel <= 24'h23_27_5F;
                10'd65: pixel <= 24'h28_5D_FF;
                10'd66: pixel <= 24'h5F_FF_23;
                10'd67: pixel <= 24'hFF_23_27;
                10'd68: pixel <= 24'h23_28_5D;
                10'd69: pixel <= 24'h28_5D_FF;
                10'd70: pixel <= 24'h5F_FF_23;
                10'd71: pixel <= 24'hFF_23_27;
                10'd72: pixel <= 24'h23_28_5D;
                10'd73: pixel <= 24'h27_5F_FF;
                10'd74: pixel <= 24'h5D_FF_23;
                10'd75: pixel <= 24'hFF_23_28;
                10'd76: pixel <= 24'h23_27_5F;
                10'd77: pixel <= 24'h28_5D_FF;
                10'd78: pixel <= 24'h5F_FF_23;
                10'd79: pixel <= 24'hFF_23_27;
                10'd80: pixel <= 24'h23_27_5F;
                10'd81: pixel <= 24'h28_5D_FF;
                10'd82: pixel <= 24'h5F_FF_23;
                10'd83: pixel <= 24'hFF_23_27;
                10'd84: pixel <= 24'h23_28_5D;
                10'd85: pixel <= 24'h27_5F_FF;
                10'd86: pixel <= 24'h7F_FF_23;
                10'd87: pixel <= 24'hFF_20_3E;
                10'd88: pixel <= 24'h38_61_AA;
                10'd89: pixel <= 24'h60_A9_FF;
                10'd90: pixel <= 24'hA9_FF_37;
                10'd91: pixel <= 24'hFF_37_60;
                10'd92: pixel <= 24'h37_60_A9;
                10'd93: pixel <= 24'h60_A9_FF;
                10'd94: pixel <= 24'hA9_FF_37;
                10'd95: pixel <= 24'hFF_37_60;
                10'd96: pixel <= 24'h37_60_A9;
                10'd97: pixel <= 24'h60_A9_FF;
                10'd98: pixel <= 24'hA9_FF_37;
                10'd99: pixel <= 24'hFF_37_60;
            endcase
            10'd25: case (x)
                10'd0: pixel <= 24'h3A_62_AB;
                10'd1: pixel <= 24'h62_AB_FF;
                10'd2: pixel <= 24'hAB_FF_3A;
                10'd3: pixel <= 24'hFF_3A_62;
                10'd4: pixel <= 24'h3A_62_AB;
                10'd5: pixel <= 24'h62_AB_FF;
                10'd6: pixel <= 24'hAB_FF_3A;
                10'd7: pixel <= 24'hFF_3A_62;
                10'd8: pixel <= 24'h3A_62_AB;
                10'd9: pixel <= 24'h62_AB_FF;
                10'd10: pixel <= 24'hAB_FF_3A;
                10'd11: pixel <= 24'hFF_3A_62;
                10'd12: pixel <= 24'h1E_41_82;
                10'd13: pixel <= 24'h27_5F_FF;
                10'd14: pixel <= 24'h5F_FF_23;
                10'd15: pixel <= 24'hFF_23_27;
                10'd16: pixel <= 24'h23_27_5F;
                10'd17: pixel <= 24'h27_5F_FF;
                10'd18: pixel <= 24'h5F_FF_23;
                10'd19: pixel <= 24'hFF_23_27;
                10'd20: pixel <= 24'h23_27_5F;
                10'd21: pixel <= 24'h27_5F_FF;
                10'd22: pixel <= 24'h5F_FF_23;
                10'd23: pixel <= 24'hFF_23_27;
                10'd24: pixel <= 24'h23_27_5F;
                10'd25: pixel <= 24'h27_5F_FF;
                10'd26: pixel <= 24'h5F_FF_23;
                10'd27: pixel <= 24'hFF_23_27;
                10'd28: pixel <= 24'h23_27_5F;
                10'd29: pixel <= 24'h27_5F_FF;
                10'd30: pixel <= 24'h5F_FF_23;
                10'd31: pixel <= 24'hFF_23_27;
                10'd32: pixel <= 24'h23_27_5F;
                10'd33: pixel <= 24'h27_5F_FF;
                10'd34: pixel <= 24'h5F_FF_23;
                10'd35: pixel <= 24'hFF_23_27;
                10'd36: pixel <= 24'h23_27_5F;
                10'd37: pixel <= 24'h27_5F_FF;
                10'd38: pixel <= 24'h5F_FF_23;
                10'd39: pixel <= 24'hFF_23_27;
                10'd40: pixel <= 24'h23_27_5F;
                10'd41: pixel <= 24'h27_5F_FF;
                10'd42: pixel <= 24'h5F_FF_23;
                10'd43: pixel <= 24'hFF_23_27;
                10'd44: pixel <= 24'h23_27_5F;
                10'd45: pixel <= 24'h27_5F_FF;
                10'd46: pixel <= 24'h5F_FF_23;
                10'd47: pixel <= 24'hFF_23_27;
                10'd48: pixel <= 24'h23_27_5F;
                10'd49: pixel <= 24'h27_5F_FF;
                10'd50: pixel <= 24'h5F_FF_23;
                10'd51: pixel <= 24'hFF_23_27;
                10'd52: pixel <= 24'h23_27_5F;
                10'd53: pixel <= 24'h3E_7F_FF;
                10'd54: pixel <= 24'hAB_FF_20;
                10'd55: pixel <= 24'hFF_3A_62;
                10'd56: pixel <= 24'h3A_62_AB;
                10'd57: pixel <= 24'h62_AB_FF;
                10'd58: pixel <= 24'hAB_FF_3A;
                10'd59: pixel <= 24'hFF_3A_62;
                10'd60: pixel <= 24'h3A_62_AB;
                10'd61: pixel <= 24'h62_AB_FF;
                10'd62: pixel <= 24'hAB_FF_3A;
                10'd63: pixel <= 24'hFF_3A_62;
                10'd64: pixel <= 24'h3A_62_AB;
                10'd65: pixel <= 24'h62_AB_FF;
                10'd66: pixel <= 24'hAB_FF_3A;
                10'd67: pixel <= 24'hFF_3A_62;
                10'd68: pixel <= 24'h3A_62_AB;
                10'd69: pixel <= 24'h62_AB_FF;
                10'd70: pixel <= 24'hAB_FF_3A;
                10'd71: pixel <= 24'hFF_3A_62;
                10'd72: pixel <= 24'h3A_62_AB;
                10'd73: pixel <= 24'h62_AB_FF;
                10'd74: pixel <= 24'hAB_FF_3A;
                10'd75: pixel <= 24'hFF_3A_62;
                10'd76: pixel <= 24'h3A_62_AB;
                10'd77: pixel <= 24'h62_AB_FF;
                10'd78: pixel <= 24'hAB_FF_3A;
                10'd79: pixel <= 24'hFF_3A_62;
                10'd80: pixel <= 24'h3A_62_AB;
                10'd81: pixel <= 24'h62_AB_FF;
                10'd82: pixel <= 24'hAB_FF_3A;
                10'd83: pixel <= 24'hFF_3A_62;
                10'd84: pixel <= 24'h3A_62_AB;
                10'd85: pixel <= 24'h62_AB_FF;
                10'd86: pixel <= 24'hAB_FF_3A;
                10'd87: pixel <= 24'hFF_3A_62;
                10'd88: pixel <= 24'h3A_62_AB;
                10'd89: pixel <= 24'h62_AB_FF;
                10'd90: pixel <= 24'hAB_FF_3A;
                10'd91: pixel <= 24'hFF_3A_62;
                10'd92: pixel <= 24'h3A_62_AB;
                10'd93: pixel <= 24'h62_AB_FF;
                10'd94: pixel <= 24'hAB_FF_3A;
                10'd95: pixel <= 24'hFF_3A_62;
                10'd96: pixel <= 24'h3A_62_AB;
                10'd97: pixel <= 24'h62_AB_FF;
                10'd98: pixel <= 24'h82_FF_3A;
                10'd99: pixel <= 24'hFF_22_40;
            endcase
            10'd26: case (x)
                10'd0: pixel <= 24'h24_28_60;
                10'd1: pixel <= 24'h28_60_FF;
                10'd2: pixel <= 24'h60_FF_24;
                10'd3: pixel <= 24'hFF_24_28;
                10'd4: pixel <= 24'h24_28_60;
                10'd5: pixel <= 24'h28_61_FF;
                10'd6: pixel <= 24'h60_FF_24;
                10'd7: pixel <= 24'hFF_24_28;
                10'd8: pixel <= 24'h24_28_60;
                10'd9: pixel <= 24'h28_60_FF;
                10'd10: pixel <= 24'h61_FF_24;
                10'd11: pixel <= 24'hFF_24_28;
                10'd12: pixel <= 24'h24_28_60;
                10'd13: pixel <= 24'h28_60_FF;
                10'd14: pixel <= 24'h60_FF_24;
                10'd15: pixel <= 24'hFF_24_28;
                10'd16: pixel <= 24'h24_28_60;
                10'd17: pixel <= 24'h28_61_FF;
                10'd18: pixel <= 24'h61_FF_24;
                10'd19: pixel <= 24'hFF_24_28;
                10'd20: pixel <= 24'h21_40_7E;
                10'd21: pixel <= 24'h64_AD_FF;
                10'd22: pixel <= 24'hAD_FF_3C;
                10'd23: pixel <= 24'hFF_3C_64;
                10'd24: pixel <= 24'h3B_63_AC;
                10'd25: pixel <= 24'h63_AC_FF;
                10'd26: pixel <= 24'hAC_FF_3A;
                10'd27: pixel <= 24'hFF_3B_62;
                10'd28: pixel <= 24'h3B_62_AA;
                10'd29: pixel <= 24'h63_AC_FF;
                10'd30: pixel <= 24'hAA_FF_3A;
                10'd31: pixel <= 24'hFF_3A_63;
                10'd32: pixel <= 24'h3A_63_AC;
                10'd33: pixel <= 24'h63_AB_FF;
                10'd34: pixel <= 24'hAB_FF_3A;
                10'd35: pixel <= 24'hFF_3A_63;
                10'd36: pixel <= 24'h3A_63_AC;
                10'd37: pixel <= 24'h63_AA_FF;
                10'd38: pixel <= 24'hAC_FF_3A;
                10'd39: pixel <= 24'hFF_3A_63;
                10'd40: pixel <= 24'h3A_63_AA;
                10'd41: pixel <= 24'h63_AC_FF;
                10'd42: pixel <= 24'hAA_FF_3A;
                10'd43: pixel <= 24'hFF_3A_63;
                10'd44: pixel <= 24'h3A_63_AC;
                10'd45: pixel <= 24'h63_AC_FF;
                10'd46: pixel <= 24'hAA_FF_3A;
                10'd47: pixel <= 24'hFF_3A_63;
                10'd48: pixel <= 24'h3A_63_AC;
                10'd49: pixel <= 24'h63_AA_FF;
                10'd50: pixel <= 24'hAC_FF_3A;
                10'd51: pixel <= 24'hFF_3A_63;
                10'd52: pixel <= 24'h3A_63_AA;
                10'd53: pixel <= 24'h63_AC_FF;
                10'd54: pixel <= 24'hAB_FF_3A;
                10'd55: pixel <= 24'hFF_3A_63;
                10'd56: pixel <= 24'h3A_63_AB;
                10'd57: pixel <= 24'h63_AC_FF;
                10'd58: pixel <= 24'hAA_FF_3A;
                10'd59: pixel <= 24'hFF_3A_63;
                10'd60: pixel <= 24'h3A_63_AC;
                10'd61: pixel <= 24'h63_AA_FF;
                10'd62: pixel <= 24'hAC_FF_3A;
                10'd63: pixel <= 24'hFF_3A_63;
                10'd64: pixel <= 24'h3A_63_AA;
                10'd65: pixel <= 24'h40_80_FF;
                10'd66: pixel <= 24'h81_FF_20;
                10'd67: pixel <= 24'hFF_24_40;
                10'd68: pixel <= 24'h3A_62_AB;
                10'd69: pixel <= 24'h62_AB_FF;
                10'd70: pixel <= 24'hAB_FF_3A;
                10'd71: pixel <= 24'hFF_3A_62;
                10'd72: pixel <= 24'h3A_62_AB;
                10'd73: pixel <= 24'h62_AB_FF;
                10'd74: pixel <= 24'hAB_FF_3A;
                10'd75: pixel <= 24'hFF_3A_62;
                10'd76: pixel <= 24'h3A_62_AB;
                10'd77: pixel <= 24'h62_AB_FF;
                10'd78: pixel <= 24'hAB_FF_3A;
                10'd79: pixel <= 24'hFF_3A_62;
                10'd80: pixel <= 24'h3A_62_AB;
                10'd81: pixel <= 24'h62_AB_FF;
                10'd82: pixel <= 24'hAB_FF_3A;
                10'd83: pixel <= 24'hFF_3A_62;
                10'd84: pixel <= 24'h3A_62_AB;
                10'd85: pixel <= 24'h62_AB_FF;
                10'd86: pixel <= 24'hAB_FF_3A;
                10'd87: pixel <= 24'hFF_3A_62;
                10'd88: pixel <= 24'h3A_62_AB;
                10'd89: pixel <= 24'h62_AB_FF;
                10'd90: pixel <= 24'hAB_FF_3A;
                10'd91: pixel <= 24'hFF_3A_62;
                10'd92: pixel <= 24'h3A_62_AB;
                10'd93: pixel <= 24'h62_AB_FF;
                10'd94: pixel <= 24'hAB_FF_3A;
                10'd95: pixel <= 24'hFF_3A_62;
                10'd96: pixel <= 24'h3A_62_AB;
                10'd97: pixel <= 24'h62_AB_FF;
                10'd98: pixel <= 24'hAB_FF_3A;
                10'd99: pixel <= 24'hFF_3A_62;
            endcase
            10'd27: case (x)
                10'd0: pixel <= 24'h24_42_85;
                10'd1: pixel <= 24'h43_86_F7;
                10'd2: pixel <= 24'h88_F7_24;
                10'd3: pixel <= 24'hF7_26_42;
                10'd4: pixel <= 24'h24_43_86;
                10'd5: pixel <= 24'h42_88_F7;
                10'd6: pixel <= 24'h86_F7_26;
                10'd7: pixel <= 24'hF7_24_43;
                10'd8: pixel <= 24'h26_42_88;
                10'd9: pixel <= 24'h42_85_F7;
                10'd10: pixel <= 24'h85_F7_24;
                10'd11: pixel <= 24'hF7_24_42;
                10'd12: pixel <= 24'h24_42_85;
                10'd13: pixel <= 24'h41_84_F7;
                10'd14: pixel <= 24'h86_F7_23;
                10'd15: pixel <= 24'hF7_24_41;
                10'd16: pixel <= 24'h23_41_84;
                10'd17: pixel <= 24'h41_86_F7;
                10'd18: pixel <= 24'h84_F7_24;
                10'd19: pixel <= 24'hF7_23_41;
                10'd20: pixel <= 24'h24_41_86;
                10'd21: pixel <= 24'h41_84_F7;
                10'd22: pixel <= 24'h84_F7_23;
                10'd23: pixel <= 24'hF7_23_41;
                10'd24: pixel <= 24'h24_41_86;
                10'd25: pixel <= 24'h41_84_F7;
                10'd26: pixel <= 24'h86_F7_23;
                10'd27: pixel <= 24'hF7_24_41;
                10'd28: pixel <= 24'h23_41_84;
                10'd29: pixel <= 24'h41_86_F7;
                10'd30: pixel <= 24'h82_F7_24;
                10'd31: pixel <= 24'hF7_23_42;
                10'd32: pixel <= 24'h24_42_80;
                10'd33: pixel <= 24'h41_81_F7;
                10'd34: pixel <= 24'hAB_FF_22;
                10'd35: pixel <= 24'hFF_38_62;
                10'd36: pixel <= 24'h38_62_A9;
                10'd37: pixel <= 24'h62_AB_FF;
                10'd38: pixel <= 24'hAB_FF_38;
                10'd39: pixel <= 24'hFF_38_62;
                10'd40: pixel <= 24'h38_62_A9;
                10'd41: pixel <= 24'h62_AB_FF;
                10'd42: pixel <= 24'hA9_FF_38;
                10'd43: pixel <= 24'hFF_38_62;
                10'd44: pixel <= 24'h38_62_AB;
                10'd45: pixel <= 24'h62_A9_FF;
                10'd46: pixel <= 24'hAB_FF_38;
                10'd47: pixel <= 24'hFF_3A_61;
                10'd48: pixel <= 24'h38_62_AB;
                10'd49: pixel <= 24'h62_AB_FF;
                10'd50: pixel <= 24'hAB_FF_38;
                10'd51: pixel <= 24'hFF_38_62;
                10'd52: pixel <= 24'h38_62_A9;
                10'd53: pixel <= 24'h62_AB_FF;
                10'd54: pixel <= 24'hA9_FF_38;
                10'd55: pixel <= 24'hFF_38_62;
                10'd56: pixel <= 24'h3A_61_AB;
                10'd57: pixel <= 24'h62_A9_FF;
                10'd58: pixel <= 24'hAB_FF_38;
                10'd59: pixel <= 24'hFF_38_62;
                10'd60: pixel <= 24'h38_62_AB;
                10'd61: pixel <= 24'h62_A9_FF;
                10'd62: pixel <= 24'hAB_FF_38;
                10'd63: pixel <= 24'hFF_38_62;
                10'd64: pixel <= 24'h38_62_A9;
                10'd65: pixel <= 24'h62_AB_FF;
                10'd66: pixel <= 24'hA9_FF_38;
                10'd67: pixel <= 24'hFF_38_62;
                10'd68: pixel <= 24'h3A_61_AB;
                10'd69: pixel <= 24'h62_AB_FF;
                10'd70: pixel <= 24'hAB_FF_38;
                10'd71: pixel <= 24'hFF_38_62;
                10'd72: pixel <= 24'h38_62_AB;
                10'd73: pixel <= 24'h62_A9_FF;
                10'd74: pixel <= 24'hAD_FF_38;
                10'd75: pixel <= 24'hFF_3A_62;
                10'd76: pixel <= 24'h3C_64_AD;
                10'd77: pixel <= 24'h64_AD_FF;
                10'd78: pixel <= 24'h83_FF_3C;
                10'd79: pixel <= 24'hFF_20_41;
                10'd80: pixel <= 24'h24_29_60;
                10'd81: pixel <= 24'h29_62_FF;
                10'd82: pixel <= 24'h60_FF_24;
                10'd83: pixel <= 24'hFF_24_28;
                10'd84: pixel <= 24'h24_28_60;
                10'd85: pixel <= 24'h28_60_FF;
                10'd86: pixel <= 24'h61_FF_24;
                10'd87: pixel <= 24'hFF_24_28;
                10'd88: pixel <= 24'h24_28_60;
                10'd89: pixel <= 24'h28_60_FF;
                10'd90: pixel <= 24'h60_FF_24;
                10'd91: pixel <= 24'hFF_24_28;
                10'd92: pixel <= 24'h24_28_60;
                10'd93: pixel <= 24'h28_61_FF;
                10'd94: pixel <= 24'h60_FF_24;
                10'd95: pixel <= 24'hFF_24_28;
                10'd96: pixel <= 24'h24_28_60;
                10'd97: pixel <= 24'h28_60_FF;
                10'd98: pixel <= 24'h61_FF_24;
                10'd99: pixel <= 24'hFF_24_28;
            endcase
            10'd28: case (x)
                10'd0: pixel <= 24'h25_43_84;
                10'd1: pixel <= 24'h42_86_F7;
                10'd2: pixel <= 24'h85_F7_25;
                10'd3: pixel <= 24'hF7_24_41;
                10'd4: pixel <= 24'h25_43_86;
                10'd5: pixel <= 24'h43_86_F7;
                10'd6: pixel <= 24'h86_F7_25;
                10'd7: pixel <= 24'hF7_25_42;
                10'd8: pixel <= 24'h25_41_88;
                10'd9: pixel <= 24'h42_86_F7;
                10'd10: pixel <= 24'h88_F7_25;
                10'd11: pixel <= 24'hF7_25_41;
                10'd12: pixel <= 24'h25_42_86;
                10'd13: pixel <= 24'h41_88_F7;
                10'd14: pixel <= 24'h84_F7_25;
                10'd15: pixel <= 24'hF7_24_41;
                10'd16: pixel <= 24'h25_42_86;
                10'd17: pixel <= 24'h41_88_F7;
                10'd18: pixel <= 24'h86_F7_25;
                10'd19: pixel <= 24'hF7_25_42;
                10'd20: pixel <= 24'h25_41_88;
                10'd21: pixel <= 24'h42_86_F7;
                10'd22: pixel <= 24'h88_F7_25;
                10'd23: pixel <= 24'hF7_25_41;
                10'd24: pixel <= 24'h24_41_84;
                10'd25: pixel <= 24'h42_86_F7;
                10'd26: pixel <= 24'h86_F7_25;
                10'd27: pixel <= 24'hF7_25_42;
                10'd28: pixel <= 24'h25_42_86;
                10'd29: pixel <= 24'h41_88_F7;
                10'd30: pixel <= 24'h86_F7_25;
                10'd31: pixel <= 24'hF7_25_42;
                10'd32: pixel <= 24'h25_41_88;
                10'd33: pixel <= 24'h42_86_F7;
                10'd34: pixel <= 24'h88_F7_25;
                10'd35: pixel <= 24'hF7_25_41;
                10'd36: pixel <= 24'h24_41_84;
                10'd37: pixel <= 24'h42_86_F7;
                10'd38: pixel <= 24'h88_F7_25;
                10'd39: pixel <= 24'hF7_25_41;
                10'd40: pixel <= 24'h23_44_84;
                10'd41: pixel <= 24'h64_AB_F8;
                10'd42: pixel <= 24'hAD_FF_40;
                10'd43: pixel <= 24'hFF_3C_64;
                10'd44: pixel <= 24'h3C_64_AD;
                10'd45: pixel <= 24'h41_85_FF;
                10'd46: pixel <= 24'h63_FF_21;
                10'd47: pixel <= 24'hFF_25_29;
                10'd48: pixel <= 24'h25_29_63;
                10'd49: pixel <= 24'h2A_61_FF;
                10'd50: pixel <= 24'h61_FF_25;
                10'd51: pixel <= 24'hFF_25_2A;
                10'd52: pixel <= 24'h25_2A_61;
                10'd53: pixel <= 24'h29_63_FF;
                10'd54: pixel <= 24'h61_FF_25;
                10'd55: pixel <= 24'hFF_25_2A;
                10'd56: pixel <= 24'h25_2A_61;
                10'd57: pixel <= 24'h2A_61_FF;
                10'd58: pixel <= 24'h61_FF_25;
                10'd59: pixel <= 24'hFF_25_2A;
                10'd60: pixel <= 24'h25_29_63;
                10'd61: pixel <= 24'h2A_61_FF;
                10'd62: pixel <= 24'h61_FF_25;
                10'd63: pixel <= 24'hFF_25_2A;
                10'd64: pixel <= 24'h25_2A_61;
                10'd65: pixel <= 24'h29_63_FF;
                10'd66: pixel <= 24'h61_FF_25;
                10'd67: pixel <= 24'hFF_25_2A;
                10'd68: pixel <= 24'h25_2A_61;
                10'd69: pixel <= 24'h2A_61_FF;
                10'd70: pixel <= 24'h61_FF_25;
                10'd71: pixel <= 24'hFF_25_2A;
                10'd72: pixel <= 24'h25_29_63;
                10'd73: pixel <= 24'h2A_61_FF;
                10'd74: pixel <= 24'h61_FF_25;
                10'd75: pixel <= 24'hFF_25_2A;
                10'd76: pixel <= 24'h25_2A_61;
                10'd77: pixel <= 24'h29_63_FF;
                10'd78: pixel <= 24'h61_FF_25;
                10'd79: pixel <= 24'hFF_25_2A;
                10'd80: pixel <= 24'h25_2A_61;
                10'd81: pixel <= 24'h2A_61_FF;
                10'd82: pixel <= 24'h61_FF_25;
                10'd83: pixel <= 24'hFF_25_2A;
                10'd84: pixel <= 24'h25_29_63;
                10'd85: pixel <= 24'h28_63_FF;
                10'd86: pixel <= 24'h7E_FF_27;
                10'd87: pixel <= 24'hFF_23_3F;
                10'd88: pixel <= 24'h3C_64_AD;
                10'd89: pixel <= 24'h64_AD_FF;
                10'd90: pixel <= 24'hAB_FF_3C;
                10'd91: pixel <= 24'hFF_3E_64;
                10'd92: pixel <= 24'h22_43_86;
                10'd93: pixel <= 24'h41_87_F8;
                10'd94: pixel <= 24'h86_F7_25;
                10'd95: pixel <= 24'hF7_26_42;
                10'd96: pixel <= 24'h24_43_88;
                10'd97: pixel <= 24'h43_86_F7;
                10'd98: pixel <= 24'h88_F7_24;
                10'd99: pixel <= 24'hF7_26_42;
            endcase
            10'd29: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'hAA_00_00;
                10'd7: pixel <= 24'h0C_40_55;
                10'd8: pixel <= 24'h41_66_AE;
                10'd9: pixel <= 24'h66_AE_FF;
                10'd10: pixel <= 24'hB0_FF_3D;
                10'd11: pixel <= 24'hFF_3D_65;
                10'd12: pixel <= 24'h21_41_85;
                10'd13: pixel <= 24'h29_63_FF;
                10'd14: pixel <= 24'h63_FF_25;
                10'd15: pixel <= 24'hFF_25_29;
                10'd16: pixel <= 24'h23_2A_63;
                10'd17: pixel <= 24'h29_63_FF;
                10'd18: pixel <= 24'h63_FF_25;
                10'd19: pixel <= 24'hFF_25_29;
                10'd20: pixel <= 24'h25_29_63;
                10'd21: pixel <= 24'h2A_63_FF;
                10'd22: pixel <= 24'h63_FF_23;
                10'd23: pixel <= 24'hFF_25_29;
                10'd24: pixel <= 24'h25_29_63;
                10'd25: pixel <= 24'h29_63_FF;
                10'd26: pixel <= 24'h63_FF_25;
                10'd27: pixel <= 24'hFF_25_29;
                10'd28: pixel <= 24'h23_2A_63;
                10'd29: pixel <= 24'h29_63_FF;
                10'd30: pixel <= 24'h63_FF_25;
                10'd31: pixel <= 24'hFF_25_29;
                10'd32: pixel <= 24'h25_29_63;
                10'd33: pixel <= 24'h2A_63_FF;
                10'd34: pixel <= 24'h63_FF_23;
                10'd35: pixel <= 24'hFF_25_29;
                10'd36: pixel <= 24'h25_29_63;
                10'd37: pixel <= 24'h29_63_FF;
                10'd38: pixel <= 24'h63_FF_25;
                10'd39: pixel <= 24'hFF_25_29;
                10'd40: pixel <= 24'h23_2A_63;
                10'd41: pixel <= 24'h29_63_FF;
                10'd42: pixel <= 24'h63_FF_25;
                10'd43: pixel <= 24'hFF_25_29;
                10'd44: pixel <= 24'h25_29_63;
                10'd45: pixel <= 24'h2A_63_FF;
                10'd46: pixel <= 24'h63_FF_23;
                10'd47: pixel <= 24'hFF_23_2A;
                10'd48: pixel <= 24'h25_29_63;
                10'd49: pixel <= 24'h29_63_FF;
                10'd50: pixel <= 24'h63_FF_25;
                10'd51: pixel <= 24'hFF_25_29;
                10'd52: pixel <= 24'h27_28_63;
                10'd53: pixel <= 24'h3E_7D_FF;
                10'd54: pixel <= 24'hAE_FF_21;
                10'd55: pixel <= 24'hFF_3D_66;
                10'd56: pixel <= 24'h3D_65_B0;
                10'd57: pixel <= 24'h64_AC_FF;
                10'd58: pixel <= 24'hAA_FF_40;
                10'd59: pixel <= 24'h0C_40_55;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd30: case (x)
                10'd0: pixel <= 24'h25_2B_66;
                10'd1: pixel <= 24'h2B_66_FF;
                10'd2: pixel <= 24'h66_FF_25;
                10'd3: pixel <= 24'hFF_25_2B;
                10'd4: pixel <= 24'h25_2B_66;
                10'd5: pixel <= 24'h2B_66_FF;
                10'd6: pixel <= 24'h66_FF_25;
                10'd7: pixel <= 24'hFF_25_2B;
                10'd8: pixel <= 24'h25_2B_66;
                10'd9: pixel <= 24'h2B_66_FF;
                10'd10: pixel <= 24'h66_FF_25;
                10'd11: pixel <= 24'hFF_23_2C;
                10'd12: pixel <= 24'h25_2B_66;
                10'd13: pixel <= 24'h2B_66_FF;
                10'd14: pixel <= 24'h66_FF_25;
                10'd15: pixel <= 24'hFF_25_2B;
                10'd16: pixel <= 24'h25_2B_66;
                10'd17: pixel <= 24'h2B_66_FF;
                10'd18: pixel <= 24'h66_FF_25;
                10'd19: pixel <= 24'hFF_25_2B;
                10'd20: pixel <= 24'h23_3F_7E;
                10'd21: pixel <= 24'h66_AE_FF;
                10'd22: pixel <= 24'hAE_FF_3D;
                10'd23: pixel <= 24'hFF_3D_66;
                10'd24: pixel <= 24'h40_65_AA;
                10'd25: pixel <= 24'h55_AA_FF;
                10'd26: pixel <= 24'h00_0C_40;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd31: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h55_AA_00;
                10'd74: pixel <= 24'hAC_0C_40;
                10'd75: pixel <= 24'hFF_41_66;
                10'd76: pixel <= 24'h3D_66_AE;
                10'd77: pixel <= 24'h66_AE_FF;
                10'd78: pixel <= 24'h85_FF_3D;
                10'd79: pixel <= 24'hFF_22_40;
                10'd80: pixel <= 24'h25_2B_66;
                10'd81: pixel <= 24'h2B_66_FF;
                10'd82: pixel <= 24'h66_FF_25;
                10'd83: pixel <= 24'hFF_25_2B;
                10'd84: pixel <= 24'h25_2B_66;
                10'd85: pixel <= 24'h2B_66_FF;
                10'd86: pixel <= 24'h66_FF_25;
                10'd87: pixel <= 24'hFF_25_2B;
                10'd88: pixel <= 24'h25_2B_66;
                10'd89: pixel <= 24'h2B_66_FF;
                10'd90: pixel <= 24'h66_FF_25;
                10'd91: pixel <= 24'hFF_25_2B;
                10'd92: pixel <= 24'h25_2B_66;
                10'd93: pixel <= 24'h2C_66_FF;
                10'd94: pixel <= 24'h66_FF_23;
                10'd95: pixel <= 24'hFF_25_2B;
                10'd96: pixel <= 24'h25_2B_66;
                10'd97: pixel <= 24'h2B_66_FF;
                10'd98: pixel <= 24'h66_FF_25;
                10'd99: pixel <= 24'hFF_25_2B;
            endcase
            10'd32: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h40_55_AA;
                10'd41: pixel <= 24'h67_AD_0C;
                10'd42: pixel <= 24'hB0_FF_43;
                10'd43: pixel <= 24'hFF_3E_67;
                10'd44: pixel <= 24'h3E_67_B0;
                10'd45: pixel <= 24'h3F_82_FF;
                10'd46: pixel <= 24'h67_FF_21;
                10'd47: pixel <= 24'hFF_26_2C;
                10'd48: pixel <= 24'h26_2C_67;
                10'd49: pixel <= 24'h2C_67_FF;
                10'd50: pixel <= 24'h67_FF_26;
                10'd51: pixel <= 24'hFF_26_2C;
                10'd52: pixel <= 24'h26_2C_67;
                10'd53: pixel <= 24'h2C_67_FF;
                10'd54: pixel <= 24'h67_FF_26;
                10'd55: pixel <= 24'hFF_26_2C;
                10'd56: pixel <= 24'h26_2C_67;
                10'd57: pixel <= 24'h2C_67_FF;
                10'd58: pixel <= 24'h67_FF_26;
                10'd59: pixel <= 24'hFF_26_2C;
                10'd60: pixel <= 24'h26_2C_67;
                10'd61: pixel <= 24'h2C_67_FF;
                10'd62: pixel <= 24'h67_FF_26;
                10'd63: pixel <= 24'hFF_26_2C;
                10'd64: pixel <= 24'h26_2C_67;
                10'd65: pixel <= 24'h2C_67_FF;
                10'd66: pixel <= 24'h67_FF_26;
                10'd67: pixel <= 24'hFF_26_2C;
                10'd68: pixel <= 24'h26_2C_67;
                10'd69: pixel <= 24'h2C_67_FF;
                10'd70: pixel <= 24'h67_FF_26;
                10'd71: pixel <= 24'hFF_26_2C;
                10'd72: pixel <= 24'h26_2C_67;
                10'd73: pixel <= 24'h2C_67_FF;
                10'd74: pixel <= 24'h67_FF_26;
                10'd75: pixel <= 24'hFF_26_2C;
                10'd76: pixel <= 24'h26_2C_67;
                10'd77: pixel <= 24'h2C_67_FF;
                10'd78: pixel <= 24'h67_FF_26;
                10'd79: pixel <= 24'hFF_26_2C;
                10'd80: pixel <= 24'h26_2C_67;
                10'd81: pixel <= 24'h2C_67_FF;
                10'd82: pixel <= 24'h67_FF_26;
                10'd83: pixel <= 24'hFF_26_2C;
                10'd84: pixel <= 24'h26_2C_67;
                10'd85: pixel <= 24'h2C_67_FF;
                10'd86: pixel <= 24'h7D_FF_26;
                10'd87: pixel <= 24'hFF_21_3E;
                10'd88: pixel <= 24'h3E_67_B0;
                10'd89: pixel <= 24'h67_B0_FF;
                10'd90: pixel <= 24'hAC_FF_3E;
                10'd91: pixel <= 24'hFF_41_66;
                10'd92: pixel <= 24'h40_55_AA;
                10'd93: pixel <= 24'h00_00_0C;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd33: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'hAA_00_00;
                10'd7: pixel <= 24'h0C_40_55;
                10'd8: pixel <= 24'h43_67_AF;
                10'd9: pixel <= 24'h67_B0_FF;
                10'd10: pixel <= 24'hB0_FF_3E;
                10'd11: pixel <= 24'hFF_3E_67;
                10'd12: pixel <= 24'h1F_40_82;
                10'd13: pixel <= 24'h2D_69_FF;
                10'd14: pixel <= 24'h6B_FF_27;
                10'd15: pixel <= 24'hFF_27_2D;
                10'd16: pixel <= 24'h26_2C_69;
                10'd17: pixel <= 24'h2C_69_FF;
                10'd18: pixel <= 24'h69_FF_26;
                10'd19: pixel <= 24'hFF_26_2C;
                10'd20: pixel <= 24'h26_2C_69;
                10'd21: pixel <= 24'h2C_69_FF;
                10'd22: pixel <= 24'h69_FF_26;
                10'd23: pixel <= 24'hFF_26_2C;
                10'd24: pixel <= 24'h26_2C_69;
                10'd25: pixel <= 24'h2C_69_FF;
                10'd26: pixel <= 24'h69_FF_26;
                10'd27: pixel <= 24'hFF_26_2C;
                10'd28: pixel <= 24'h26_2C_69;
                10'd29: pixel <= 24'h2C_69_FF;
                10'd30: pixel <= 24'h69_FF_26;
                10'd31: pixel <= 24'hFF_26_2C;
                10'd32: pixel <= 24'h26_2C_69;
                10'd33: pixel <= 24'h2C_69_FF;
                10'd34: pixel <= 24'h69_FF_26;
                10'd35: pixel <= 24'hFF_26_2C;
                10'd36: pixel <= 24'h26_2C_69;
                10'd37: pixel <= 24'h2C_69_FF;
                10'd38: pixel <= 24'h69_FF_26;
                10'd39: pixel <= 24'hFF_26_2C;
                10'd40: pixel <= 24'h26_2C_69;
                10'd41: pixel <= 24'h2C_69_FF;
                10'd42: pixel <= 24'h69_FF_26;
                10'd43: pixel <= 24'hFF_26_2C;
                10'd44: pixel <= 24'h26_2C_69;
                10'd45: pixel <= 24'h2C_69_FF;
                10'd46: pixel <= 24'h69_FF_26;
                10'd47: pixel <= 24'hFF_26_2C;
                10'd48: pixel <= 24'h26_2C_69;
                10'd49: pixel <= 24'h2C_69_FF;
                10'd50: pixel <= 24'h69_FF_26;
                10'd51: pixel <= 24'hFF_26_2C;
                10'd52: pixel <= 24'h26_2C_69;
                10'd53: pixel <= 24'h3E_7D_FF;
                10'd54: pixel <= 24'hB0_FF_21;
                10'd55: pixel <= 24'hFF_3E_67;
                10'd56: pixel <= 24'h3E_67_B0;
                10'd57: pixel <= 24'h66_AC_FF;
                10'd58: pixel <= 24'hAA_FF_41;
                10'd59: pixel <= 24'h0C_40_55;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd34: case (x)
                10'd0: pixel <= 24'h27_2D_6B;
                10'd1: pixel <= 24'h2D_6B_FF;
                10'd2: pixel <= 24'h6B_FF_27;
                10'd3: pixel <= 24'hFF_27_2D;
                10'd4: pixel <= 24'h27_2D_6B;
                10'd5: pixel <= 24'h2D_6B_FF;
                10'd6: pixel <= 24'h6B_FF_27;
                10'd7: pixel <= 24'hFF_27_2D;
                10'd8: pixel <= 24'h27_2D_6B;
                10'd9: pixel <= 24'h2D_6B_FF;
                10'd10: pixel <= 24'h6B_FF_27;
                10'd11: pixel <= 24'hFF_27_2D;
                10'd12: pixel <= 24'h27_2D_6B;
                10'd13: pixel <= 24'h2D_6B_FF;
                10'd14: pixel <= 24'h6B_FF_27;
                10'd15: pixel <= 24'hFF_27_2D;
                10'd16: pixel <= 24'h27_2D_6B;
                10'd17: pixel <= 24'h2D_6B_FF;
                10'd18: pixel <= 24'h6B_FF_27;
                10'd19: pixel <= 24'hFF_27_2D;
                10'd20: pixel <= 24'h21_3E_7D;
                10'd21: pixel <= 24'h68_B1_FF;
                10'd22: pixel <= 24'hB1_FF_3F;
                10'd23: pixel <= 24'hFF_3F_68;
                10'd24: pixel <= 24'h43_67_AD;
                10'd25: pixel <= 24'h55_AA_FF;
                10'd26: pixel <= 24'h00_0C_40;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd35: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h55_AA_00;
                10'd74: pixel <= 24'hAF_0C_40;
                10'd75: pixel <= 24'hFF_43_67;
                10'd76: pixel <= 24'h3F_68_B1;
                10'd77: pixel <= 24'h68_B1_FF;
                10'd78: pixel <= 24'h81_FF_3F;
                10'd79: pixel <= 24'hFF_1E_3F;
                10'd80: pixel <= 24'h27_2D_6B;
                10'd81: pixel <= 24'h2D_6B_FF;
                10'd82: pixel <= 24'h6B_FF_27;
                10'd83: pixel <= 24'hFF_27_2D;
                10'd84: pixel <= 24'h27_2D_6B;
                10'd85: pixel <= 24'h2D_6B_FF;
                10'd86: pixel <= 24'h6B_FF_27;
                10'd87: pixel <= 24'hFF_27_2D;
                10'd88: pixel <= 24'h27_2D_6B;
                10'd89: pixel <= 24'h2D_6B_FF;
                10'd90: pixel <= 24'h6B_FF_27;
                10'd91: pixel <= 24'hFF_27_2D;
                10'd92: pixel <= 24'h27_2D_6B;
                10'd93: pixel <= 24'h2D_6B_FF;
                10'd94: pixel <= 24'h6B_FF_27;
                10'd95: pixel <= 24'hFF_27_2D;
                10'd96: pixel <= 24'h27_2D_6B;
                10'd97: pixel <= 24'h2D_6B_FF;
                10'd98: pixel <= 24'h6B_FF_27;
                10'd99: pixel <= 24'hFF_27_2D;
            endcase
            10'd36: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h40_55_AA;
                10'd41: pixel <= 24'h68_B0_0C;
                10'd42: pixel <= 24'hB2_FF_44;
                10'd43: pixel <= 24'hFF_41_69;
                10'd44: pixel <= 24'h41_69_B0;
                10'd45: pixel <= 24'h3F_84_FF;
                10'd46: pixel <= 24'h6E_FF_1F;
                10'd47: pixel <= 24'hFF_28_2E;
                10'd48: pixel <= 24'h28_2E_6E;
                10'd49: pixel <= 24'h2E_6E_FF;
                10'd50: pixel <= 24'h6E_FF_28;
                10'd51: pixel <= 24'hFF_28_2E;
                10'd52: pixel <= 24'h28_2E_6E;
                10'd53: pixel <= 24'h2E_6E_FF;
                10'd54: pixel <= 24'h6E_FF_28;
                10'd55: pixel <= 24'hFF_28_2E;
                10'd56: pixel <= 24'h28_2E_6E;
                10'd57: pixel <= 24'h2E_6E_FF;
                10'd58: pixel <= 24'h6E_FF_28;
                10'd59: pixel <= 24'hFF_28_2E;
                10'd60: pixel <= 24'h28_2E_6E;
                10'd61: pixel <= 24'h2E_6E_FF;
                10'd62: pixel <= 24'h6E_FF_28;
                10'd63: pixel <= 24'hFF_28_2E;
                10'd64: pixel <= 24'h28_2E_6E;
                10'd65: pixel <= 24'h2E_6E_FF;
                10'd66: pixel <= 24'h6E_FF_28;
                10'd67: pixel <= 24'hFF_28_2E;
                10'd68: pixel <= 24'h28_2E_6E;
                10'd69: pixel <= 24'h2E_6E_FF;
                10'd70: pixel <= 24'h6E_FF_28;
                10'd71: pixel <= 24'hFF_28_2E;
                10'd72: pixel <= 24'h28_2E_6E;
                10'd73: pixel <= 24'h2E_6E_FF;
                10'd74: pixel <= 24'h6E_FF_28;
                10'd75: pixel <= 24'hFF_28_2E;
                10'd76: pixel <= 24'h28_2E_6E;
                10'd77: pixel <= 24'h2E_6E_FF;
                10'd78: pixel <= 24'h6E_FF_28;
                10'd79: pixel <= 24'hFF_28_2E;
                10'd80: pixel <= 24'h28_2E_6E;
                10'd81: pixel <= 24'h2E_6E_FF;
                10'd82: pixel <= 24'h6E_FF_28;
                10'd83: pixel <= 24'hFF_28_2E;
                10'd84: pixel <= 24'h28_2E_6E;
                10'd85: pixel <= 24'h2E_6E_FF;
                10'd86: pixel <= 24'h80_FF_28;
                10'd87: pixel <= 24'hFF_23_3F;
                10'd88: pixel <= 24'h41_69_B2;
                10'd89: pixel <= 24'h69_B2_FF;
                10'd90: pixel <= 24'hAE_FF_41;
                10'd91: pixel <= 24'hFF_44_68;
                10'd92: pixel <= 24'h40_55_AA;
                10'd93: pixel <= 24'h00_00_0C;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd37: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'hAA_00_00;
                10'd7: pixel <= 24'h0C_40_55;
                10'd8: pixel <= 24'h45_69_B1;
                10'd9: pixel <= 24'h6B_B1_FF;
                10'd10: pixel <= 24'hB3_FF_42;
                10'd11: pixel <= 24'hFF_42_6A;
                10'd12: pixel <= 24'h1E_3E_83;
                10'd13: pixel <= 24'h2F_6F_FF;
                10'd14: pixel <= 24'h71_FF_29;
                10'd15: pixel <= 24'hFF_29_2E;
                10'd16: pixel <= 24'h29_2E_71;
                10'd17: pixel <= 24'h2E_71_FF;
                10'd18: pixel <= 24'h6F_FF_29;
                10'd19: pixel <= 24'hFF_29_2F;
                10'd20: pixel <= 24'h29_2E_71;
                10'd21: pixel <= 24'h2F_71_FF;
                10'd22: pixel <= 24'h71_FF_28;
                10'd23: pixel <= 24'hFF_29_2E;
                10'd24: pixel <= 24'h29_2E_71;
                10'd25: pixel <= 24'h2E_71_FF;
                10'd26: pixel <= 24'h71_FF_29;
                10'd27: pixel <= 24'hFF_29_2E;
                10'd28: pixel <= 24'h28_30_6F;
                10'd29: pixel <= 24'h2E_71_FF;
                10'd30: pixel <= 24'h71_FF_29;
                10'd31: pixel <= 24'hFF_29_2E;
                10'd32: pixel <= 24'h29_2E_71;
                10'd33: pixel <= 24'h2F_71_FF;
                10'd34: pixel <= 24'h71_FF_28;
                10'd35: pixel <= 24'hFF_29_2E;
                10'd36: pixel <= 24'h29_2E_71;
                10'd37: pixel <= 24'h2F_6F_FF;
                10'd38: pixel <= 24'h71_FF_29;
                10'd39: pixel <= 24'hFF_29_2E;
                10'd40: pixel <= 24'h28_2F_71;
                10'd41: pixel <= 24'h2E_71_FF;
                10'd42: pixel <= 24'h71_FF_29;
                10'd43: pixel <= 24'hFF_29_2E;
                10'd44: pixel <= 24'h29_2E_71;
                10'd45: pixel <= 24'h30_6F_FF;
                10'd46: pixel <= 24'h6F_FF_28;
                10'd47: pixel <= 24'hFF_28_30;
                10'd48: pixel <= 24'h29_2E_71;
                10'd49: pixel <= 24'h2E_71_FF;
                10'd50: pixel <= 24'h71_FF_29;
                10'd51: pixel <= 24'hFF_29_2E;
                10'd52: pixel <= 24'h29_2F_6F;
                10'd53: pixel <= 24'h3D_7F_FF;
                10'd54: pixel <= 24'hB1_FF_21;
                10'd55: pixel <= 24'hFF_42_6B;
                10'd56: pixel <= 24'h42_6A_B3;
                10'd57: pixel <= 24'h69_AF_FF;
                10'd58: pixel <= 24'hAA_FF_45;
                10'd59: pixel <= 24'h0C_40_55;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd38: case (x)
                10'd0: pixel <= 24'h28_2F_71;
                10'd1: pixel <= 24'h2E_71_FF;
                10'd2: pixel <= 24'h71_FF_29;
                10'd3: pixel <= 24'hFF_29_2E;
                10'd4: pixel <= 24'h29_2F_6F;
                10'd5: pixel <= 24'h2E_71_FF;
                10'd6: pixel <= 24'h71_FF_29;
                10'd7: pixel <= 24'hFF_28_2F;
                10'd8: pixel <= 24'h29_2E_71;
                10'd9: pixel <= 24'h2E_71_FF;
                10'd10: pixel <= 24'h71_FF_29;
                10'd11: pixel <= 24'hFF_29_2E;
                10'd12: pixel <= 24'h28_30_6F;
                10'd13: pixel <= 24'h30_6F_FF;
                10'd14: pixel <= 24'h71_FF_28;
                10'd15: pixel <= 24'hFF_29_2E;
                10'd16: pixel <= 24'h29_2E_71;
                10'd17: pixel <= 24'h2E_71_FF;
                10'd18: pixel <= 24'h6F_FF_29;
                10'd19: pixel <= 24'hFF_29_2F;
                10'd20: pixel <= 24'h21_3E_7D;
                10'd21: pixel <= 24'h6B_B1_FF;
                10'd22: pixel <= 24'hB3_FF_42;
                10'd23: pixel <= 24'hFF_42_6A;
                10'd24: pixel <= 24'h45_69_AF;
                10'd25: pixel <= 24'h55_AA_FF;
                10'd26: pixel <= 24'h00_0C_40;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd39: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h55_AA_00;
                10'd74: pixel <= 24'hAF_0C_40;
                10'd75: pixel <= 24'hFF_45_69;
                10'd76: pixel <= 24'h42_6B_B1;
                10'd77: pixel <= 24'h6A_B3_FF;
                10'd78: pixel <= 24'h84_FF_42;
                10'd79: pixel <= 24'hFF_1F_3F;
                10'd80: pixel <= 24'h29_2F_6F;
                10'd81: pixel <= 24'h2E_71_FF;
                10'd82: pixel <= 24'h71_FF_29;
                10'd83: pixel <= 24'hFF_29_2E;
                10'd84: pixel <= 24'h29_2E_71;
                10'd85: pixel <= 24'h2F_6F_FF;
                10'd86: pixel <= 24'h71_FF_29;
                10'd87: pixel <= 24'hFF_29_2E;
                10'd88: pixel <= 24'h28_2F_71;
                10'd89: pixel <= 24'h2E_71_FF;
                10'd90: pixel <= 24'h71_FF_29;
                10'd91: pixel <= 24'hFF_29_2E;
                10'd92: pixel <= 24'h29_2E_71;
                10'd93: pixel <= 24'h2E_71_FF;
                10'd94: pixel <= 24'h6F_FF_29;
                10'd95: pixel <= 24'hFF_28_30;
                10'd96: pixel <= 24'h29_2E_71;
                10'd97: pixel <= 24'h2E_71_FF;
                10'd98: pixel <= 24'h71_FF_29;
                10'd99: pixel <= 24'hFF_29_2E;
            endcase
            10'd40: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h40_55_AA;
                10'd41: pixel <= 24'h69_AF_0C;
                10'd42: pixel <= 24'hB4_FF_45;
                10'd43: pixel <= 24'hFF_43_6B;
                10'd44: pixel <= 24'h43_6C_B2;
                10'd45: pixel <= 24'h3F_84_FF;
                10'd46: pixel <= 24'h70_FF_1F;
                10'd47: pixel <= 24'hFF_2A_30;
                10'd48: pixel <= 24'h2A_30_72;
                10'd49: pixel <= 24'h30_72_FF;
                10'd50: pixel <= 24'h72_FF_29;
                10'd51: pixel <= 24'hFF_29_30;
                10'd52: pixel <= 24'h29_30_72;
                10'd53: pixel <= 24'h30_72_FF;
                10'd54: pixel <= 24'h72_FF_29;
                10'd55: pixel <= 24'hFF_2A_30;
                10'd56: pixel <= 24'h29_30_72;
                10'd57: pixel <= 24'h30_72_FF;
                10'd58: pixel <= 24'h72_FF_29;
                10'd59: pixel <= 24'hFF_29_30;
                10'd60: pixel <= 24'h29_30_72;
                10'd61: pixel <= 24'h30_72_FF;
                10'd62: pixel <= 24'h72_FF_2A;
                10'd63: pixel <= 24'hFF_29_30;
                10'd64: pixel <= 24'h29_30_72;
                10'd65: pixel <= 24'h30_72_FF;
                10'd66: pixel <= 24'h72_FF_29;
                10'd67: pixel <= 24'hFF_2A_30;
                10'd68: pixel <= 24'h29_30_72;
                10'd69: pixel <= 24'h30_72_FF;
                10'd70: pixel <= 24'h72_FF_29;
                10'd71: pixel <= 24'hFF_29_30;
                10'd72: pixel <= 24'h29_30_72;
                10'd73: pixel <= 24'h30_72_FF;
                10'd74: pixel <= 24'h72_FF_2A;
                10'd75: pixel <= 24'hFF_29_30;
                10'd76: pixel <= 24'h29_30_72;
                10'd77: pixel <= 24'h30_72_FF;
                10'd78: pixel <= 24'h72_FF_29;
                10'd79: pixel <= 24'hFF_2A_30;
                10'd80: pixel <= 24'h2A_30_72;
                10'd81: pixel <= 24'h30_72_FF;
                10'd82: pixel <= 24'h72_FF_29;
                10'd83: pixel <= 24'hFF_29_30;
                10'd84: pixel <= 24'h29_30_72;
                10'd85: pixel <= 24'h30_72_FF;
                10'd86: pixel <= 24'h7E_FF_2A;
                10'd87: pixel <= 24'hFF_23_3F;
                10'd88: pixel <= 24'h43_6B_B4;
                10'd89: pixel <= 24'h6B_B4_FF;
                10'd90: pixel <= 24'hB0_FF_43;
                10'd91: pixel <= 24'hFF_46_6B;
                10'd92: pixel <= 24'h40_55_AA;
                10'd93: pixel <= 24'h00_00_0C;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd41: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'hAA_00_00;
                10'd7: pixel <= 24'h0C_40_55;
                10'd8: pixel <= 24'h46_6B_B0;
                10'd9: pixel <= 24'h6C_B2_FF;
                10'd10: pixel <= 24'hB2_FF_43;
                10'd11: pixel <= 24'hFF_43_6C;
                10'd12: pixel <= 24'h1E_3E_85;
                10'd13: pixel <= 24'h30_72_FF;
                10'd14: pixel <= 24'h74_FF_2A;
                10'd15: pixel <= 24'hFF_2A_2F;
                10'd16: pixel <= 24'h29_30_74;
                10'd17: pixel <= 24'h30_74_FF;
                10'd18: pixel <= 24'h74_FF_29;
                10'd19: pixel <= 24'hFF_29_30;
                10'd20: pixel <= 24'h29_30_74;
                10'd21: pixel <= 24'h30_74_FF;
                10'd22: pixel <= 24'h74_FF_29;
                10'd23: pixel <= 24'hFF_29_30;
                10'd24: pixel <= 24'h29_30_74;
                10'd25: pixel <= 24'h30_74_FF;
                10'd26: pixel <= 24'h74_FF_29;
                10'd27: pixel <= 24'hFF_29_30;
                10'd28: pixel <= 24'h29_30_74;
                10'd29: pixel <= 24'h30_74_FF;
                10'd30: pixel <= 24'h74_FF_29;
                10'd31: pixel <= 24'hFF_29_30;
                10'd32: pixel <= 24'h29_30_74;
                10'd33: pixel <= 24'h30_74_FF;
                10'd34: pixel <= 24'h74_FF_29;
                10'd35: pixel <= 24'hFF_29_30;
                10'd36: pixel <= 24'h29_30_74;
                10'd37: pixel <= 24'h30_74_FF;
                10'd38: pixel <= 24'h74_FF_29;
                10'd39: pixel <= 24'hFF_29_30;
                10'd40: pixel <= 24'h29_30_74;
                10'd41: pixel <= 24'h30_74_FF;
                10'd42: pixel <= 24'h74_FF_29;
                10'd43: pixel <= 24'hFF_29_30;
                10'd44: pixel <= 24'h29_30_74;
                10'd45: pixel <= 24'h30_74_FF;
                10'd46: pixel <= 24'h74_FF_29;
                10'd47: pixel <= 24'hFF_29_30;
                10'd48: pixel <= 24'h29_30_74;
                10'd49: pixel <= 24'h30_74_FF;
                10'd50: pixel <= 24'h74_FF_29;
                10'd51: pixel <= 24'hFF_29_30;
                10'd52: pixel <= 24'h2A_30_72;
                10'd53: pixel <= 24'h3F_7E_FF;
                10'd54: pixel <= 24'hB2_FF_23;
                10'd55: pixel <= 24'hFF_43_6C;
                10'd56: pixel <= 24'h43_6C_B2;
                10'd57: pixel <= 24'h6B_AE_FF;
                10'd58: pixel <= 24'hAA_FF_46;
                10'd59: pixel <= 24'h0C_40_55;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd42: case (x)
                10'd0: pixel <= 24'h2A_31_75;
                10'd1: pixel <= 24'h31_75_FF;
                10'd2: pixel <= 24'h75_FF_2A;
                10'd3: pixel <= 24'hFF_2A_31;
                10'd4: pixel <= 24'h2A_31_75;
                10'd5: pixel <= 24'h31_75_FF;
                10'd6: pixel <= 24'h75_FF_2A;
                10'd7: pixel <= 24'hFF_2A_31;
                10'd8: pixel <= 24'h2A_31_75;
                10'd9: pixel <= 24'h31_75_FF;
                10'd10: pixel <= 24'h75_FF_2A;
                10'd11: pixel <= 24'hFF_2A_31;
                10'd12: pixel <= 24'h2A_31_75;
                10'd13: pixel <= 24'h31_75_FF;
                10'd14: pixel <= 24'h75_FF_2A;
                10'd15: pixel <= 24'hFF_2A_31;
                10'd16: pixel <= 24'h2A_31_75;
                10'd17: pixel <= 24'h31_75_FF;
                10'd18: pixel <= 24'h75_FF_2A;
                10'd19: pixel <= 24'hFF_2A_31;
                10'd20: pixel <= 24'h23_3F_7E;
                10'd21: pixel <= 24'h6D_B3_FF;
                10'd22: pixel <= 24'hB3_FF_44;
                10'd23: pixel <= 24'hFF_44_6D;
                10'd24: pixel <= 24'h47_6C_AF;
                10'd25: pixel <= 24'h55_AA_FF;
                10'd26: pixel <= 24'h00_0C_40;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd43: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h55_AA_00;
                10'd74: pixel <= 24'hB0_0C_40;
                10'd75: pixel <= 24'hFF_46_6B;
                10'd76: pixel <= 24'h44_6D_B3;
                10'd77: pixel <= 24'h6D_B3_FF;
                10'd78: pixel <= 24'h86_FF_44;
                10'd79: pixel <= 24'hFF_1F_3F;
                10'd80: pixel <= 24'h2A_31_73;
                10'd81: pixel <= 24'h31_75_FF;
                10'd82: pixel <= 24'h75_FF_2A;
                10'd83: pixel <= 24'hFF_2A_31;
                10'd84: pixel <= 24'h2A_31_75;
                10'd85: pixel <= 24'h31_75_FF;
                10'd86: pixel <= 24'h75_FF_2A;
                10'd87: pixel <= 24'hFF_2A_31;
                10'd88: pixel <= 24'h2A_31_75;
                10'd89: pixel <= 24'h31_75_FF;
                10'd90: pixel <= 24'h75_FF_2A;
                10'd91: pixel <= 24'hFF_2A_31;
                10'd92: pixel <= 24'h2A_31_75;
                10'd93: pixel <= 24'h31_75_FF;
                10'd94: pixel <= 24'h75_FF_2A;
                10'd95: pixel <= 24'hFF_2A_31;
                10'd96: pixel <= 24'h2A_31_75;
                10'd97: pixel <= 24'h31_75_FF;
                10'd98: pixel <= 24'h75_FF_2A;
                10'd99: pixel <= 24'hFF_2A_31;
            endcase
            10'd44: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h40_55_AA;
                10'd41: pixel <= 24'h6D_B3_0C;
                10'd42: pixel <= 24'hB5_FF_48;
                10'd43: pixel <= 24'hFF_45_6E;
                10'd44: pixel <= 24'h45_6E_B5;
                10'd45: pixel <= 24'h3F_84_FF;
                10'd46: pixel <= 24'h76_FF_1F;
                10'd47: pixel <= 24'hFF_2B_32;
                10'd48: pixel <= 24'h2B_32_78;
                10'd49: pixel <= 24'h32_78_FF;
                10'd50: pixel <= 24'h78_FF_2B;
                10'd51: pixel <= 24'hFF_2B_32;
                10'd52: pixel <= 24'h2B_32_78;
                10'd53: pixel <= 24'h32_78_FF;
                10'd54: pixel <= 24'h78_FF_2B;
                10'd55: pixel <= 24'hFF_2B_32;
                10'd56: pixel <= 24'h2B_32_78;
                10'd57: pixel <= 24'h32_78_FF;
                10'd58: pixel <= 24'h78_FF_2B;
                10'd59: pixel <= 24'hFF_2B_32;
                10'd60: pixel <= 24'h2B_32_78;
                10'd61: pixel <= 24'h32_78_FF;
                10'd62: pixel <= 24'h78_FF_2B;
                10'd63: pixel <= 24'hFF_2B_32;
                10'd64: pixel <= 24'h2B_32_78;
                10'd65: pixel <= 24'h32_78_FF;
                10'd66: pixel <= 24'h78_FF_2B;
                10'd67: pixel <= 24'hFF_2B_32;
                10'd68: pixel <= 24'h2B_32_78;
                10'd69: pixel <= 24'h32_78_FF;
                10'd70: pixel <= 24'h78_FF_2B;
                10'd71: pixel <= 24'hFF_2B_32;
                10'd72: pixel <= 24'h2B_32_78;
                10'd73: pixel <= 24'h32_78_FF;
                10'd74: pixel <= 24'h78_FF_2B;
                10'd75: pixel <= 24'hFF_2B_32;
                10'd76: pixel <= 24'h2B_32_78;
                10'd77: pixel <= 24'h32_78_FF;
                10'd78: pixel <= 24'h78_FF_2B;
                10'd79: pixel <= 24'hFF_2B_32;
                10'd80: pixel <= 24'h2B_32_78;
                10'd81: pixel <= 24'h32_78_FF;
                10'd82: pixel <= 24'h78_FF_2B;
                10'd83: pixel <= 24'hFF_2B_32;
                10'd84: pixel <= 24'h2B_32_78;
                10'd85: pixel <= 24'h32_76_FF;
                10'd86: pixel <= 24'h7D_FF_2B;
                10'd87: pixel <= 24'hFF_21_3E;
                10'd88: pixel <= 24'h44_6D_B3;
                10'd89: pixel <= 24'h6D_B3_FF;
                10'd90: pixel <= 24'hAF_FF_44;
                10'd91: pixel <= 24'hFF_47_6C;
                10'd92: pixel <= 24'h40_55_AA;
                10'd93: pixel <= 24'h00_00_0C;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd45: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'hAA_00_00;
                10'd7: pixel <= 24'h0C_40_55;
                10'd8: pixel <= 24'h48_6D_B3;
                10'd9: pixel <= 24'h6E_B5_FF;
                10'd10: pixel <= 24'hB3_FF_45;
                10'd11: pixel <= 24'hFF_45_6F;
                10'd12: pixel <= 24'h1F_3F_84;
                10'd13: pixel <= 24'h33_78_FF;
                10'd14: pixel <= 24'h7A_FF_2C;
                10'd15: pixel <= 24'hFF_2C_33;
                10'd16: pixel <= 24'h2C_33_7A;
                10'd17: pixel <= 24'h33_7A_FF;
                10'd18: pixel <= 24'h7A_FF_2C;
                10'd19: pixel <= 24'hFF_2C_33;
                10'd20: pixel <= 24'h2C_33_7A;
                10'd21: pixel <= 24'h33_7A_FF;
                10'd22: pixel <= 24'h7C_FF_2C;
                10'd23: pixel <= 24'hFF_2C_33;
                10'd24: pixel <= 24'h2C_33_7A;
                10'd25: pixel <= 24'h33_7A_FF;
                10'd26: pixel <= 24'h7A_FF_2C;
                10'd27: pixel <= 24'hFF_2C_33;
                10'd28: pixel <= 24'h2C_33_7A;
                10'd29: pixel <= 24'h33_7C_FF;
                10'd30: pixel <= 24'h7A_FF_2C;
                10'd31: pixel <= 24'hFF_2C_33;
                10'd32: pixel <= 24'h2C_33_7A;
                10'd33: pixel <= 24'h33_7A_FF;
                10'd34: pixel <= 24'h7C_FF_2C;
                10'd35: pixel <= 24'hFF_2C_33;
                10'd36: pixel <= 24'h2C_33_7C;
                10'd37: pixel <= 24'h33_7A_FF;
                10'd38: pixel <= 24'h7A_FF_2C;
                10'd39: pixel <= 24'hFF_2C_33;
                10'd40: pixel <= 24'h2C_33_7A;
                10'd41: pixel <= 24'h33_7C_FF;
                10'd42: pixel <= 24'h7A_FF_2C;
                10'd43: pixel <= 24'hFF_2C_33;
                10'd44: pixel <= 24'h2C_33_7A;
                10'd45: pixel <= 24'h33_7A_FF;
                10'd46: pixel <= 24'h7A_FF_2C;
                10'd47: pixel <= 24'hFF_2C_33;
                10'd48: pixel <= 24'h2C_33_7C;
                10'd49: pixel <= 24'h33_7A_FF;
                10'd50: pixel <= 24'h7A_FF_2C;
                10'd51: pixel <= 24'hFF_2C_33;
                10'd52: pixel <= 24'h2C_33_7A;
                10'd53: pixel <= 24'h3F_7E_FF;
                10'd54: pixel <= 24'hB5_FF_23;
                10'd55: pixel <= 24'hFF_45_6E;
                10'd56: pixel <= 24'h45_6E_B5;
                10'd57: pixel <= 24'h6D_B1_FF;
                10'd58: pixel <= 24'hAA_FF_48;
                10'd59: pixel <= 24'h0C_40_55;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd46: case (x)
                10'd0: pixel <= 24'h2C_33_7C;
                10'd1: pixel <= 24'h33_7C_FF;
                10'd2: pixel <= 24'h7C_FF_2C;
                10'd3: pixel <= 24'hFF_2C_33;
                10'd4: pixel <= 24'h2C_33_7C;
                10'd5: pixel <= 24'h33_7C_FF;
                10'd6: pixel <= 24'h7C_FF_2C;
                10'd7: pixel <= 24'hFF_2C_33;
                10'd8: pixel <= 24'h2C_33_7C;
                10'd9: pixel <= 24'h33_7C_FF;
                10'd10: pixel <= 24'h7C_FF_2C;
                10'd11: pixel <= 24'hFF_2C_33;
                10'd12: pixel <= 24'h2C_33_7C;
                10'd13: pixel <= 24'h33_7C_FF;
                10'd14: pixel <= 24'h7C_FF_2C;
                10'd15: pixel <= 24'hFF_2C_33;
                10'd16: pixel <= 24'h2C_33_7C;
                10'd17: pixel <= 24'h33_7C_FF;
                10'd18: pixel <= 24'h7A_FF_2C;
                10'd19: pixel <= 24'hFF_2C_33;
                10'd20: pixel <= 24'h22_3E_7D;
                10'd21: pixel <= 24'h6F_B6_FF;
                10'd22: pixel <= 24'hB6_FF_46;
                10'd23: pixel <= 24'hFF_46_6F;
                10'd24: pixel <= 24'h4A_6E_B2;
                10'd25: pixel <= 24'h55_AA_FF;
                10'd26: pixel <= 24'h00_0C_40;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd47: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h55_AA_00;
                10'd74: pixel <= 24'hB6_0C_40;
                10'd75: pixel <= 24'hFF_4A_6E;
                10'd76: pixel <= 24'h46_6F_B6;
                10'd77: pixel <= 24'h6F_B6_FF;
                10'd78: pixel <= 24'h86_FF_46;
                10'd79: pixel <= 24'hFF_1F_3F;
                10'd80: pixel <= 24'h2C_33_7A;
                10'd81: pixel <= 24'h33_7C_FF;
                10'd82: pixel <= 24'h7C_FF_2C;
                10'd83: pixel <= 24'hFF_2C_33;
                10'd84: pixel <= 24'h2C_33_7C;
                10'd85: pixel <= 24'h33_7C_FF;
                10'd86: pixel <= 24'h7C_FF_2C;
                10'd87: pixel <= 24'hFF_2C_33;
                10'd88: pixel <= 24'h2C_33_7C;
                10'd89: pixel <= 24'h33_7C_FF;
                10'd90: pixel <= 24'h7C_FF_2C;
                10'd91: pixel <= 24'hFF_2C_33;
                10'd92: pixel <= 24'h2C_33_7C;
                10'd93: pixel <= 24'h33_7C_FF;
                10'd94: pixel <= 24'h7C_FF_2C;
                10'd95: pixel <= 24'hFF_2C_33;
                10'd96: pixel <= 24'h2C_33_7C;
                10'd97: pixel <= 24'h33_7C_FF;
                10'd98: pixel <= 24'h7C_FF_2C;
                10'd99: pixel <= 24'hFF_2C_33;
            endcase
            10'd48: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h40_55_AA;
                10'd41: pixel <= 24'h6F_B7_0C;
                10'd42: pixel <= 24'hB5_FF_4B;
                10'd43: pixel <= 24'hFF_48_71;
                10'd44: pixel <= 24'h48_71_B5;
                10'd45: pixel <= 24'h3F_84_FF;
                10'd46: pixel <= 24'h7A_FF_1F;
                10'd47: pixel <= 24'hFF_2C_33;
                10'd48: pixel <= 24'h2C_33_7C;
                10'd49: pixel <= 24'h33_7C_FF;
                10'd50: pixel <= 24'h7C_FF_2C;
                10'd51: pixel <= 24'hFF_2C_33;
                10'd52: pixel <= 24'h2C_33_7C;
                10'd53: pixel <= 24'h33_7C_FF;
                10'd54: pixel <= 24'h7C_FF_2C;
                10'd55: pixel <= 24'hFF_2C_33;
                10'd56: pixel <= 24'h2C_33_7C;
                10'd57: pixel <= 24'h33_7C_FF;
                10'd58: pixel <= 24'h7C_FF_2C;
                10'd59: pixel <= 24'hFF_2C_33;
                10'd60: pixel <= 24'h2C_33_7C;
                10'd61: pixel <= 24'h33_7C_FF;
                10'd62: pixel <= 24'h7C_FF_2C;
                10'd63: pixel <= 24'hFF_2C_33;
                10'd64: pixel <= 24'h2C_33_7C;
                10'd65: pixel <= 24'h33_7C_FF;
                10'd66: pixel <= 24'h7C_FF_2C;
                10'd67: pixel <= 24'hFF_2C_33;
                10'd68: pixel <= 24'h2C_33_7C;
                10'd69: pixel <= 24'h33_7C_FF;
                10'd70: pixel <= 24'h7C_FF_2C;
                10'd71: pixel <= 24'hFF_2C_33;
                10'd72: pixel <= 24'h2C_33_7C;
                10'd73: pixel <= 24'h33_7C_FF;
                10'd74: pixel <= 24'h7C_FF_2C;
                10'd75: pixel <= 24'hFF_2C_33;
                10'd76: pixel <= 24'h2C_33_7C;
                10'd77: pixel <= 24'h33_7C_FF;
                10'd78: pixel <= 24'h7C_FF_2C;
                10'd79: pixel <= 24'hFF_2C_33;
                10'd80: pixel <= 24'h2C_33_7C;
                10'd81: pixel <= 24'h33_7C_FF;
                10'd82: pixel <= 24'h7C_FF_2C;
                10'd83: pixel <= 24'hFF_2C_33;
                10'd84: pixel <= 24'h2C_33_7C;
                10'd85: pixel <= 24'h33_7A_FF;
                10'd86: pixel <= 24'h82_FF_2C;
                10'd87: pixel <= 24'hFF_26_42;
                10'd88: pixel <= 24'h48_70_B7;
                10'd89: pixel <= 24'h71_B5_FF;
                10'd90: pixel <= 24'hB3_FF_48;
                10'd91: pixel <= 24'hFF_4B_70;
                10'd92: pixel <= 24'h40_55_AA;
                10'd93: pixel <= 24'h00_00_0C;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd49: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'hAA_00_00;
                10'd7: pixel <= 24'h0C_40_55;
                10'd8: pixel <= 24'h4B_6F_B7;
                10'd9: pixel <= 24'h72_B6_FF;
                10'd10: pixel <= 24'hB7_FF_49;
                10'd11: pixel <= 24'hFF_49_72;
                10'd12: pixel <= 24'h1F_40_82;
                10'd13: pixel <= 24'h33_7B_FF;
                10'd14: pixel <= 24'h7C_FF_2C;
                10'd15: pixel <= 24'hFF_2C_33;
                10'd16: pixel <= 24'h2C_33_7C;
                10'd17: pixel <= 24'h33_7D_FF;
                10'd18: pixel <= 24'h7C_FF_2C;
                10'd19: pixel <= 24'hFF_2C_33;
                10'd20: pixel <= 24'h2C_33_7D;
                10'd21: pixel <= 24'h33_7C_FF;
                10'd22: pixel <= 24'h7D_FF_2C;
                10'd23: pixel <= 24'hFF_2C_33;
                10'd24: pixel <= 24'h2C_33_7C;
                10'd25: pixel <= 24'h33_7C_FF;
                10'd26: pixel <= 24'h7D_FF_2C;
                10'd27: pixel <= 24'hFF_2C_33;
                10'd28: pixel <= 24'h2C_33_7C;
                10'd29: pixel <= 24'h33_7D_FF;
                10'd30: pixel <= 24'h7C_FF_2C;
                10'd31: pixel <= 24'hFF_2C_33;
                10'd32: pixel <= 24'h2C_33_7D;
                10'd33: pixel <= 24'h33_7C_FF;
                10'd34: pixel <= 24'h7D_FF_2C;
                10'd35: pixel <= 24'hFF_2C_33;
                10'd36: pixel <= 24'h2C_33_7D;
                10'd37: pixel <= 24'h33_7C_FF;
                10'd38: pixel <= 24'h7D_FF_2C;
                10'd39: pixel <= 24'hFF_2C_33;
                10'd40: pixel <= 24'h2C_33_7C;
                10'd41: pixel <= 24'h33_7D_FF;
                10'd42: pixel <= 24'h7C_FF_2C;
                10'd43: pixel <= 24'hFF_2C_33;
                10'd44: pixel <= 24'h2C_33_7D;
                10'd45: pixel <= 24'h33_7C_FF;
                10'd46: pixel <= 24'h7C_FF_2C;
                10'd47: pixel <= 24'hFF_2C_33;
                10'd48: pixel <= 24'h2C_33_7D;
                10'd49: pixel <= 24'h33_7C_FF;
                10'd50: pixel <= 24'h7D_FF_2C;
                10'd51: pixel <= 24'hFF_2C_33;
                10'd52: pixel <= 24'h2C_33_7B;
                10'd53: pixel <= 24'h42_82_FF;
                10'd54: pixel <= 24'hB8_FF_26;
                10'd55: pixel <= 24'hFF_49_72;
                10'd56: pixel <= 24'h49_72_B7;
                10'd57: pixel <= 24'h71_B4_FF;
                10'd58: pixel <= 24'hAA_FF_4C;
                10'd59: pixel <= 24'h0C_40_55;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd50: case (x)
                10'd0: pixel <= 24'h2C_33_7C;
                10'd1: pixel <= 24'h32_7E_FF;
                10'd2: pixel <= 24'h7E_FF_2C;
                10'd3: pixel <= 24'hFF_2C_32;
                10'd4: pixel <= 24'h2C_33_7C;
                10'd5: pixel <= 24'h32_7E_FF;
                10'd6: pixel <= 24'h7C_FF_2C;
                10'd7: pixel <= 24'hFF_2C_33;
                10'd8: pixel <= 24'h2C_32_7E;
                10'd9: pixel <= 24'h33_7C_FF;
                10'd10: pixel <= 24'h7E_FF_2C;
                10'd11: pixel <= 24'hFF_2C_32;
                10'd12: pixel <= 24'h2C_33_7C;
                10'd13: pixel <= 24'h33_7C_FF;
                10'd14: pixel <= 24'h7E_FF_2C;
                10'd15: pixel <= 24'hFF_2C_32;
                10'd16: pixel <= 24'h2C_33_7C;
                10'd17: pixel <= 24'h32_7E_FF;
                10'd18: pixel <= 24'h7C_FF_2C;
                10'd19: pixel <= 24'hFF_2C_33;
                10'd20: pixel <= 24'h25_41_81;
                10'd21: pixel <= 24'h71_B8_FF;
                10'd22: pixel <= 24'hB8_FF_4A;
                10'd23: pixel <= 24'hFF_49_72;
                10'd24: pixel <= 24'h4C_71_B4;
                10'd25: pixel <= 24'h55_AA_FF;
                10'd26: pixel <= 24'h00_0C_40;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd51: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h55_AA_00;
                10'd74: pixel <= 24'hB7_0C_40;
                10'd75: pixel <= 24'hFF_4C_70;
                10'd76: pixel <= 24'h4A_71_B6;
                10'd77: pixel <= 24'h72_B8_FF;
                10'd78: pixel <= 24'h82_FF_49;
                10'd79: pixel <= 24'hFF_1F_40;
                10'd80: pixel <= 24'h2C_33_7C;
                10'd81: pixel <= 24'h33_7C_FF;
                10'd82: pixel <= 24'h7C_FF_2C;
                10'd83: pixel <= 24'hFF_2C_33;
                10'd84: pixel <= 24'h2C_32_7E;
                10'd85: pixel <= 24'h33_7C_FF;
                10'd86: pixel <= 24'h7E_FF_2C;
                10'd87: pixel <= 24'hFF_2C_32;
                10'd88: pixel <= 24'h2C_33_7C;
                10'd89: pixel <= 24'h32_7E_FF;
                10'd90: pixel <= 24'h7C_FF_2C;
                10'd91: pixel <= 24'hFF_2C_33;
                10'd92: pixel <= 24'h2C_33_7C;
                10'd93: pixel <= 24'h32_7E_FF;
                10'd94: pixel <= 24'h7C_FF_2C;
                10'd95: pixel <= 24'hFF_2C_33;
                10'd96: pixel <= 24'h2C_32_7E;
                10'd97: pixel <= 24'h33_7C_FF;
                10'd98: pixel <= 24'h7E_FF_2C;
                10'd99: pixel <= 24'hFF_2C_32;
            endcase
            10'd52: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h40_55_AA;
                10'd41: pixel <= 24'h70_B6_0C;
                10'd42: pixel <= 24'hB7_FF_4C;
                10'd43: pixel <= 24'hFF_4C_72;
                10'd44: pixel <= 24'h4C_72_B7;
                10'd45: pixel <= 24'h40_82_FF;
                10'd46: pixel <= 24'h7E_FF_1F;
                10'd47: pixel <= 24'hFF_2C_32;
                10'd48: pixel <= 24'h2C_32_7E;
                10'd49: pixel <= 24'h32_7E_FF;
                10'd50: pixel <= 24'h7E_FF_2C;
                10'd51: pixel <= 24'hFF_2C_32;
                10'd52: pixel <= 24'h2C_32_7E;
                10'd53: pixel <= 24'h32_7E_FF;
                10'd54: pixel <= 24'h7E_FF_2C;
                10'd55: pixel <= 24'hFF_2C_32;
                10'd56: pixel <= 24'h2C_32_7E;
                10'd57: pixel <= 24'h32_7E_FF;
                10'd58: pixel <= 24'h7E_FF_2C;
                10'd59: pixel <= 24'hFF_2C_32;
                10'd60: pixel <= 24'h2C_32_7E;
                10'd61: pixel <= 24'h32_7E_FF;
                10'd62: pixel <= 24'h7E_FF_2C;
                10'd63: pixel <= 24'hFF_2C_32;
                10'd64: pixel <= 24'h2C_32_7E;
                10'd65: pixel <= 24'h32_7E_FF;
                10'd66: pixel <= 24'h7E_FF_2C;
                10'd67: pixel <= 24'hFF_2C_32;
                10'd68: pixel <= 24'h2C_32_7E;
                10'd69: pixel <= 24'h32_7E_FF;
                10'd70: pixel <= 24'h7E_FF_2C;
                10'd71: pixel <= 24'hFF_2C_32;
                10'd72: pixel <= 24'h2C_32_7E;
                10'd73: pixel <= 24'h32_7E_FF;
                10'd74: pixel <= 24'h7E_FF_2C;
                10'd75: pixel <= 24'hFF_2C_32;
                10'd76: pixel <= 24'h2C_32_7E;
                10'd77: pixel <= 24'h32_7E_FF;
                10'd78: pixel <= 24'h7E_FF_2C;
                10'd79: pixel <= 24'hFF_2C_32;
                10'd80: pixel <= 24'h2C_32_7E;
                10'd81: pixel <= 24'h32_7E_FF;
                10'd82: pixel <= 24'h7E_FF_2C;
                10'd83: pixel <= 24'hFF_2C_32;
                10'd84: pixel <= 24'h2C_32_7E;
                10'd85: pixel <= 24'h32_7C_FF;
                10'd86: pixel <= 24'h83_FF_2E;
                10'd87: pixel <= 24'hFF_25_41;
                10'd88: pixel <= 24'h4C_72_B7;
                10'd89: pixel <= 24'h72_B7_FF;
                10'd90: pixel <= 24'hB5_FF_4C;
                10'd91: pixel <= 24'hFF_4D_72;
                10'd92: pixel <= 24'h40_55_AA;
                10'd93: pixel <= 24'h00_00_0C;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd53: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'hAA_00_00;
                10'd7: pixel <= 24'h0C_40_55;
                10'd8: pixel <= 24'h4D_72_B7;
                10'd9: pixel <= 24'h72_B7_FF;
                10'd10: pixel <= 24'hB7_FF_4C;
                10'd11: pixel <= 24'hFF_4C_72;
                10'd12: pixel <= 24'h1F_40_82;
                10'd13: pixel <= 24'h32_7E_FF;
                10'd14: pixel <= 24'h7E_FF_2C;
                10'd15: pixel <= 24'hFF_2C_32;
                10'd16: pixel <= 24'h2E_31_7E;
                10'd17: pixel <= 24'h32_7E_FF;
                10'd18: pixel <= 24'h7E_FF_2C;
                10'd19: pixel <= 24'hFF_2E_31;
                10'd20: pixel <= 24'h2C_32_7E;
                10'd21: pixel <= 24'h31_7E_FF;
                10'd22: pixel <= 24'h7E_FF_2E;
                10'd23: pixel <= 24'hFF_2C_32;
                10'd24: pixel <= 24'h2E_31_7E;
                10'd25: pixel <= 24'h31_7E_FF;
                10'd26: pixel <= 24'h7E_FF_2E;
                10'd27: pixel <= 24'hFF_2C_32;
                10'd28: pixel <= 24'h2E_31_7E;
                10'd29: pixel <= 24'h32_7E_FF;
                10'd30: pixel <= 24'h7E_FF_2C;
                10'd31: pixel <= 24'hFF_2E_31;
                10'd32: pixel <= 24'h2C_32_7E;
                10'd33: pixel <= 24'h31_7E_FF;
                10'd34: pixel <= 24'h7E_FF_2E;
                10'd35: pixel <= 24'hFF_2C_32;
                10'd36: pixel <= 24'h2C_32_7E;
                10'd37: pixel <= 24'h31_7E_FF;
                10'd38: pixel <= 24'h7E_FF_2E;
                10'd39: pixel <= 24'hFF_2C_32;
                10'd40: pixel <= 24'h2E_31_7E;
                10'd41: pixel <= 24'h32_7E_FF;
                10'd42: pixel <= 24'h7E_FF_2C;
                10'd43: pixel <= 24'hFF_2E_31;
                10'd44: pixel <= 24'h2C_32_7E;
                10'd45: pixel <= 24'h31_7E_FF;
                10'd46: pixel <= 24'h7E_FF_2E;
                10'd47: pixel <= 24'hFF_2E_31;
                10'd48: pixel <= 24'h2C_32_7E;
                10'd49: pixel <= 24'h31_7E_FF;
                10'd50: pixel <= 24'h7E_FF_2E;
                10'd51: pixel <= 24'hFF_2C_32;
                10'd52: pixel <= 24'h2E_32_7C;
                10'd53: pixel <= 24'h42_84_FF;
                10'd54: pixel <= 24'hB7_FF_26;
                10'd55: pixel <= 24'hFF_4C_72;
                10'd56: pixel <= 24'h4C_72_B7;
                10'd57: pixel <= 24'h72_B5_FF;
                10'd58: pixel <= 24'hAA_FF_4D;
                10'd59: pixel <= 24'h0C_40_55;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd54: case (x)
                10'd0: pixel <= 24'h2C_32_7E;
                10'd1: pixel <= 24'h32_7E_FF;
                10'd2: pixel <= 24'h7E_FF_2C;
                10'd3: pixel <= 24'hFF_2C_32;
                10'd4: pixel <= 24'h2C_32_7E;
                10'd5: pixel <= 24'h32_7E_FF;
                10'd6: pixel <= 24'h7E_FF_2C;
                10'd7: pixel <= 24'hFF_2C_32;
                10'd8: pixel <= 24'h2C_32_7E;
                10'd9: pixel <= 24'h32_7E_FF;
                10'd10: pixel <= 24'h7E_FF_2C;
                10'd11: pixel <= 24'hFF_2C_32;
                10'd12: pixel <= 24'h2C_32_7E;
                10'd13: pixel <= 24'h32_7E_FF;
                10'd14: pixel <= 24'h7E_FF_2C;
                10'd15: pixel <= 24'hFF_2C_32;
                10'd16: pixel <= 24'h2C_32_7E;
                10'd17: pixel <= 24'h32_7E_FF;
                10'd18: pixel <= 24'h7D_FF_2C;
                10'd19: pixel <= 24'hFF_2E_31;
                10'd20: pixel <= 24'h26_42_84;
                10'd21: pixel <= 24'h74_B8_FF;
                10'd22: pixel <= 24'hB8_FF_4D;
                10'd23: pixel <= 24'hFF_4D_74;
                10'd24: pixel <= 24'h4E_73_B6;
                10'd25: pixel <= 24'h55_AA_FF;
                10'd26: pixel <= 24'h00_0C_40;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd55: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h55_AA_00;
                10'd74: pixel <= 24'hB8_0C_40;
                10'd75: pixel <= 24'hFF_50_72;
                10'd76: pixel <= 24'h4D_74_B8;
                10'd77: pixel <= 24'h74_B8_FF;
                10'd78: pixel <= 24'h84_FF_4D;
                10'd79: pixel <= 24'hFF_1F_3F;
                10'd80: pixel <= 24'h2C_32_7E;
                10'd81: pixel <= 24'h32_7E_FF;
                10'd82: pixel <= 24'h7E_FF_2C;
                10'd83: pixel <= 24'hFF_2C_32;
                10'd84: pixel <= 24'h2C_32_7E;
                10'd85: pixel <= 24'h32_7E_FF;
                10'd86: pixel <= 24'h7E_FF_2C;
                10'd87: pixel <= 24'hFF_2C_32;
                10'd88: pixel <= 24'h2C_32_7E;
                10'd89: pixel <= 24'h32_7E_FF;
                10'd90: pixel <= 24'h7E_FF_2C;
                10'd91: pixel <= 24'hFF_2C_32;
                10'd92: pixel <= 24'h2C_32_7E;
                10'd93: pixel <= 24'h32_7E_FF;
                10'd94: pixel <= 24'h7E_FF_2C;
                10'd95: pixel <= 24'hFF_2C_32;
                10'd96: pixel <= 24'h2C_32_7E;
                10'd97: pixel <= 24'h32_7E_FF;
                10'd98: pixel <= 24'h7E_FF_2C;
                10'd99: pixel <= 24'hFF_2C_32;
            endcase
            10'd56: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h40_55_AA;
                10'd41: pixel <= 24'h74_BB_0C;
                10'd42: pixel <= 24'hBA_FF_52;
                10'd43: pixel <= 24'hFF_4E_75;
                10'd44: pixel <= 24'h4E_75_BA;
                10'd45: pixel <= 24'h3F_84_FF;
                10'd46: pixel <= 24'h7E_FF_1F;
                10'd47: pixel <= 24'hFF_2C_32;
                10'd48: pixel <= 24'h2C_32_7E;
                10'd49: pixel <= 24'h32_80_FF;
                10'd50: pixel <= 24'h7E_FF_2C;
                10'd51: pixel <= 24'hFF_2C_32;
                10'd52: pixel <= 24'h2C_32_80;
                10'd53: pixel <= 24'h32_7E_FF;
                10'd54: pixel <= 24'h80_FF_2C;
                10'd55: pixel <= 24'hFF_2C_32;
                10'd56: pixel <= 24'h2C_32_7E;
                10'd57: pixel <= 24'h32_80_FF;
                10'd58: pixel <= 24'h80_FF_2C;
                10'd59: pixel <= 24'hFF_2C_32;
                10'd60: pixel <= 24'h2C_32_7E;
                10'd61: pixel <= 24'h32_80_FF;
                10'd62: pixel <= 24'h7E_FF_2C;
                10'd63: pixel <= 24'hFF_2C_32;
                10'd64: pixel <= 24'h2C_32_80;
                10'd65: pixel <= 24'h32_7E_FF;
                10'd66: pixel <= 24'h80_FF_2C;
                10'd67: pixel <= 24'hFF_2C_32;
                10'd68: pixel <= 24'h2C_32_7E;
                10'd69: pixel <= 24'h32_7E_FF;
                10'd70: pixel <= 24'h80_FF_2C;
                10'd71: pixel <= 24'hFF_2C_32;
                10'd72: pixel <= 24'h2C_32_7E;
                10'd73: pixel <= 24'h32_80_FF;
                10'd74: pixel <= 24'h7E_FF_2C;
                10'd75: pixel <= 24'hFF_2C_32;
                10'd76: pixel <= 24'h2C_32_80;
                10'd77: pixel <= 24'h32_7E_FF;
                10'd78: pixel <= 24'h80_FF_2C;
                10'd79: pixel <= 24'hFF_2C_32;
                10'd80: pixel <= 24'h2C_32_80;
                10'd81: pixel <= 24'h32_7E_FF;
                10'd82: pixel <= 24'h80_FF_2C;
                10'd83: pixel <= 24'hFF_2C_32;
                10'd84: pixel <= 24'h2C_32_7E;
                10'd85: pixel <= 24'h32_7E_FF;
                10'd86: pixel <= 24'h84_FF_2C;
                10'd87: pixel <= 24'hFF_26_42;
                10'd88: pixel <= 24'h4E_75_BA;
                10'd89: pixel <= 24'h75_BA_FF;
                10'd90: pixel <= 24'hB8_FF_4E;
                10'd91: pixel <= 24'hFF_4F_74;
                10'd92: pixel <= 24'h40_55_AA;
                10'd93: pixel <= 24'h00_00_0C;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd57: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'hAA_00_00;
                10'd7: pixel <= 24'h0C_40_55;
                10'd8: pixel <= 24'h52_74_BB;
                10'd9: pixel <= 24'h75_BA_FF;
                10'd10: pixel <= 24'hBA_FF_4E;
                10'd11: pixel <= 24'hFF_4E_75;
                10'd12: pixel <= 24'h1F_3F_84;
                10'd13: pixel <= 24'h32_80_FF;
                10'd14: pixel <= 24'h80_FF_2C;
                10'd15: pixel <= 24'hFF_2C_32;
                10'd16: pixel <= 24'h2C_32_80;
                10'd17: pixel <= 24'h32_80_FF;
                10'd18: pixel <= 24'h80_FF_2C;
                10'd19: pixel <= 24'hFF_2C_32;
                10'd20: pixel <= 24'h2C_32_80;
                10'd21: pixel <= 24'h32_80_FF;
                10'd22: pixel <= 24'h80_FF_2C;
                10'd23: pixel <= 24'hFF_2C_32;
                10'd24: pixel <= 24'h2C_32_80;
                10'd25: pixel <= 24'h32_80_FF;
                10'd26: pixel <= 24'h80_FF_2C;
                10'd27: pixel <= 24'hFF_2C_32;
                10'd28: pixel <= 24'h2C_32_80;
                10'd29: pixel <= 24'h32_80_FF;
                10'd30: pixel <= 24'h80_FF_2C;
                10'd31: pixel <= 24'hFF_2C_32;
                10'd32: pixel <= 24'h2C_32_80;
                10'd33: pixel <= 24'h32_80_FF;
                10'd34: pixel <= 24'h80_FF_2C;
                10'd35: pixel <= 24'hFF_2C_32;
                10'd36: pixel <= 24'h2C_32_80;
                10'd37: pixel <= 24'h32_80_FF;
                10'd38: pixel <= 24'h80_FF_2C;
                10'd39: pixel <= 24'hFF_2C_32;
                10'd40: pixel <= 24'h2C_32_80;
                10'd41: pixel <= 24'h32_80_FF;
                10'd42: pixel <= 24'h80_FF_2C;
                10'd43: pixel <= 24'hFF_2C_32;
                10'd44: pixel <= 24'h2C_32_80;
                10'd45: pixel <= 24'h32_80_FF;
                10'd46: pixel <= 24'h80_FF_2C;
                10'd47: pixel <= 24'hFF_2C_32;
                10'd48: pixel <= 24'h2C_32_80;
                10'd49: pixel <= 24'h32_80_FF;
                10'd50: pixel <= 24'h80_FF_2C;
                10'd51: pixel <= 24'hFF_2C_32;
                10'd52: pixel <= 24'h2E_31_80;
                10'd53: pixel <= 24'h42_82_FF;
                10'd54: pixel <= 24'hBA_FF_26;
                10'd55: pixel <= 24'hFF_4E_75;
                10'd56: pixel <= 24'h4E_75_BA;
                10'd57: pixel <= 24'h74_B8_FF;
                10'd58: pixel <= 24'hAA_FF_4F;
                10'd59: pixel <= 24'h0C_40_55;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd58: case (x)
                10'd0: pixel <= 24'h2C_32_80;
                10'd1: pixel <= 24'h32_80_FF;
                10'd2: pixel <= 24'h80_FF_2C;
                10'd3: pixel <= 24'hFF_2C_32;
                10'd4: pixel <= 24'h2C_32_80;
                10'd5: pixel <= 24'h32_80_FF;
                10'd6: pixel <= 24'h80_FF_2C;
                10'd7: pixel <= 24'hFF_2C_32;
                10'd8: pixel <= 24'h2C_32_80;
                10'd9: pixel <= 24'h32_80_FF;
                10'd10: pixel <= 24'h80_FF_2C;
                10'd11: pixel <= 24'hFF_2C_32;
                10'd12: pixel <= 24'h2C_32_80;
                10'd13: pixel <= 24'h32_80_FF;
                10'd14: pixel <= 24'h80_FF_2C;
                10'd15: pixel <= 24'hFF_2C_32;
                10'd16: pixel <= 24'h2C_32_80;
                10'd17: pixel <= 24'h32_80_FF;
                10'd18: pixel <= 24'h80_FF_2C;
                10'd19: pixel <= 24'hFF_2C_32;
                10'd20: pixel <= 24'h25_41_81;
                10'd21: pixel <= 24'h76_B9_FF;
                10'd22: pixel <= 24'hB9_FF_4F;
                10'd23: pixel <= 24'hFF_4F_76;
                10'd24: pixel <= 24'h52_75_B7;
                10'd25: pixel <= 24'h55_AA_FF;
                10'd26: pixel <= 24'h00_0C_40;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd59: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h55_AA_00;
                10'd74: pixel <= 24'hB9_0C_40;
                10'd75: pixel <= 24'hFF_52_75;
                10'd76: pixel <= 24'h4F_76_B9;
                10'd77: pixel <= 24'h76_B9_FF;
                10'd78: pixel <= 24'h84_FF_4F;
                10'd79: pixel <= 24'hFF_1F_3F;
                10'd80: pixel <= 24'h2C_32_80;
                10'd81: pixel <= 24'h32_80_FF;
                10'd82: pixel <= 24'h80_FF_2C;
                10'd83: pixel <= 24'hFF_2C_32;
                10'd84: pixel <= 24'h2C_32_80;
                10'd85: pixel <= 24'h32_80_FF;
                10'd86: pixel <= 24'h80_FF_2C;
                10'd87: pixel <= 24'hFF_2C_32;
                10'd88: pixel <= 24'h2C_32_80;
                10'd89: pixel <= 24'h32_80_FF;
                10'd90: pixel <= 24'h80_FF_2C;
                10'd91: pixel <= 24'hFF_2C_32;
                10'd92: pixel <= 24'h2C_32_80;
                10'd93: pixel <= 24'h32_80_FF;
                10'd94: pixel <= 24'h80_FF_2C;
                10'd95: pixel <= 24'hFF_2C_32;
                10'd96: pixel <= 24'h2C_32_80;
                10'd97: pixel <= 24'h32_80_FF;
                10'd98: pixel <= 24'h80_FF_2C;
                10'd99: pixel <= 24'hFF_2C_32;
            endcase
            10'd60: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h40_55_AA;
                10'd41: pixel <= 24'h77_BB_0C;
                10'd42: pixel <= 24'hBA_FF_55;
                10'd43: pixel <= 24'hFF_50_77;
                10'd44: pixel <= 24'h50_77_BA;
                10'd45: pixel <= 24'h3F_84_FF;
                10'd46: pixel <= 24'h80_FF_1F;
                10'd47: pixel <= 24'hFF_2C_32;
                10'd48: pixel <= 24'h2C_32_80;
                10'd49: pixel <= 24'h32_80_FF;
                10'd50: pixel <= 24'h80_FF_2C;
                10'd51: pixel <= 24'hFF_2C_32;
                10'd52: pixel <= 24'h2C_32_80;
                10'd53: pixel <= 24'h32_80_FF;
                10'd54: pixel <= 24'h80_FF_2C;
                10'd55: pixel <= 24'hFF_2C_32;
                10'd56: pixel <= 24'h2C_32_80;
                10'd57: pixel <= 24'h32_80_FF;
                10'd58: pixel <= 24'h80_FF_2C;
                10'd59: pixel <= 24'hFF_2C_32;
                10'd60: pixel <= 24'h2C_32_80;
                10'd61: pixel <= 24'h32_80_FF;
                10'd62: pixel <= 24'h80_FF_2C;
                10'd63: pixel <= 24'hFF_2C_32;
                10'd64: pixel <= 24'h2C_32_80;
                10'd65: pixel <= 24'h32_80_FF;
                10'd66: pixel <= 24'h80_FF_2C;
                10'd67: pixel <= 24'hFF_2C_32;
                10'd68: pixel <= 24'h2C_32_80;
                10'd69: pixel <= 24'h32_80_FF;
                10'd70: pixel <= 24'h80_FF_2C;
                10'd71: pixel <= 24'hFF_2C_32;
                10'd72: pixel <= 24'h2C_32_80;
                10'd73: pixel <= 24'h32_80_FF;
                10'd74: pixel <= 24'h80_FF_2C;
                10'd75: pixel <= 24'hFF_2C_32;
                10'd76: pixel <= 24'h2C_32_80;
                10'd77: pixel <= 24'h32_80_FF;
                10'd78: pixel <= 24'h80_FF_2C;
                10'd79: pixel <= 24'hFF_2C_32;
                10'd80: pixel <= 24'h2C_32_80;
                10'd81: pixel <= 24'h32_80_FF;
                10'd82: pixel <= 24'h80_FF_2C;
                10'd83: pixel <= 24'hFF_2C_32;
                10'd84: pixel <= 24'h2C_32_80;
                10'd85: pixel <= 24'h32_80_FF;
                10'd86: pixel <= 24'h81_FF_2C;
                10'd87: pixel <= 24'hFF_25_41;
                10'd88: pixel <= 24'h50_77_BA;
                10'd89: pixel <= 24'h77_BA_FF;
                10'd90: pixel <= 24'hB8_FF_50;
                10'd91: pixel <= 24'hFF_52_77;
                10'd92: pixel <= 24'h40_55_AA;
                10'd93: pixel <= 24'h00_00_0C;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd61: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'hAA_00_00;
                10'd7: pixel <= 24'h0C_40_55;
                10'd8: pixel <= 24'h55_77_BB;
                10'd9: pixel <= 24'h77_BA_FF;
                10'd10: pixel <= 24'hBA_FF_50;
                10'd11: pixel <= 24'hFF_50_77;
                10'd12: pixel <= 24'h1F_3F_84;
                10'd13: pixel <= 24'h33_80_FF;
                10'd14: pixel <= 24'h80_FF_2B;
                10'd15: pixel <= 24'hFF_2B_33;
                10'd16: pixel <= 24'h2B_33_80;
                10'd17: pixel <= 24'h33_80_FF;
                10'd18: pixel <= 24'h80_FF_2B;
                10'd19: pixel <= 24'hFF_2B_33;
                10'd20: pixel <= 24'h2B_33_80;
                10'd21: pixel <= 24'h33_80_FF;
                10'd22: pixel <= 24'h80_FF_2B;
                10'd23: pixel <= 24'hFF_2B_33;
                10'd24: pixel <= 24'h2B_33_80;
                10'd25: pixel <= 24'h33_80_FF;
                10'd26: pixel <= 24'h80_FF_2B;
                10'd27: pixel <= 24'hFF_2B_33;
                10'd28: pixel <= 24'h2B_33_80;
                10'd29: pixel <= 24'h33_80_FF;
                10'd30: pixel <= 24'h80_FF_2B;
                10'd31: pixel <= 24'hFF_2B_33;
                10'd32: pixel <= 24'h2B_33_80;
                10'd33: pixel <= 24'h33_80_FF;
                10'd34: pixel <= 24'h80_FF_2B;
                10'd35: pixel <= 24'hFF_2B_33;
                10'd36: pixel <= 24'h2B_33_80;
                10'd37: pixel <= 24'h33_80_FF;
                10'd38: pixel <= 24'h80_FF_2B;
                10'd39: pixel <= 24'hFF_2B_33;
                10'd40: pixel <= 24'h2B_33_80;
                10'd41: pixel <= 24'h33_80_FF;
                10'd42: pixel <= 24'h80_FF_2B;
                10'd43: pixel <= 24'hFF_2B_33;
                10'd44: pixel <= 24'h2B_33_80;
                10'd45: pixel <= 24'h33_80_FF;
                10'd46: pixel <= 24'h80_FF_2B;
                10'd47: pixel <= 24'hFF_2C_32;
                10'd48: pixel <= 24'h2C_32_80;
                10'd49: pixel <= 24'h32_80_FF;
                10'd50: pixel <= 24'h80_FF_2C;
                10'd51: pixel <= 24'hFF_2E_31;
                10'd52: pixel <= 24'h2C_32_80;
                10'd53: pixel <= 24'h41_81_FF;
                10'd54: pixel <= 24'hBA_FF_25;
                10'd55: pixel <= 24'hFF_50_77;
                10'd56: pixel <= 24'h50_77_BA;
                10'd57: pixel <= 24'h77_B8_FF;
                10'd58: pixel <= 24'hAA_FF_52;
                10'd59: pixel <= 24'h0C_40_55;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd62: case (x)
                10'd0: pixel <= 24'h28_38_84;
                10'd1: pixel <= 24'h37_84_FF;
                10'd2: pixel <= 24'h84_FF_29;
                10'd3: pixel <= 24'hFF_29_36;
                10'd4: pixel <= 24'h29_36_84;
                10'd5: pixel <= 24'h36_84_FF;
                10'd6: pixel <= 24'h84_FF_29;
                10'd7: pixel <= 24'hFF_29_36;
                10'd8: pixel <= 24'h29_36_84;
                10'd9: pixel <= 24'h35_83_FF;
                10'd10: pixel <= 24'h83_FF_28;
                10'd11: pixel <= 24'hFF_28_35;
                10'd12: pixel <= 24'h28_35_81;
                10'd13: pixel <= 24'h34_7E_FF;
                10'd14: pixel <= 24'h81_FF_26;
                10'd15: pixel <= 24'hFF_29_35;
                10'd16: pixel <= 24'h2A_36_7F;
                10'd17: pixel <= 24'h35_81_FF;
                10'd18: pixel <= 24'h7F_FF_2A;
                10'd19: pixel <= 24'hFF_2C_34;
                10'd20: pixel <= 24'h25_41_83;
                10'd21: pixel <= 24'h79_BB_FF;
                10'd22: pixel <= 24'hBB_FF_51;
                10'd23: pixel <= 24'hFF_51_79;
                10'd24: pixel <= 24'h53_78_B9;
                10'd25: pixel <= 24'h55_AA_FF;
                10'd26: pixel <= 24'h00_0C_40;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd63: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h55_AA_00;
                10'd74: pixel <= 24'hBC_0C_40;
                10'd75: pixel <= 24'hFF_56_78;
                10'd76: pixel <= 24'h51_79_BB;
                10'd77: pixel <= 24'h79_BB_FF;
                10'd78: pixel <= 24'h87_FF_51;
                10'd79: pixel <= 24'hFF_21_40;
                10'd80: pixel <= 24'h29_35_83;
                10'd81: pixel <= 24'h36_83_FF;
                10'd82: pixel <= 24'h83_FF_28;
                10'd83: pixel <= 24'hFF_28_35;
                10'd84: pixel <= 24'h26_36_83;
                10'd85: pixel <= 24'h36_82_FF;
                10'd86: pixel <= 24'h82_FF_25;
                10'd87: pixel <= 24'hFF_27_35;
                10'd88: pixel <= 24'h28_35_83;
                10'd89: pixel <= 24'h35_83_FF;
                10'd90: pixel <= 24'h83_FF_28;
                10'd91: pixel <= 24'hFF_27_35;
                10'd92: pixel <= 24'h28_36_83;
                10'd93: pixel <= 24'h35_83_FF;
                10'd94: pixel <= 24'h82_FF_28;
                10'd95: pixel <= 24'hFF_27_34;
                10'd96: pixel <= 24'h27_34_82;
                10'd97: pixel <= 24'h35_83_FF;
                10'd98: pixel <= 24'h85_FF_28;
                10'd99: pixel <= 24'hFF_2B_38;
            endcase
            10'd64: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h40_55_AA;
                10'd41: pixel <= 24'h78_BC_0C;
                10'd42: pixel <= 24'hBC_FF_56;
                10'd43: pixel <= 24'hFF_52_7A;
                10'd44: pixel <= 24'h52_7A_BC;
                10'd45: pixel <= 24'h75_B8_FF;
                10'd46: pixel <= 24'hB7_FF_50;
                10'd47: pixel <= 24'hFF_4F_74;
                10'd48: pixel <= 24'h52_74_B8;
                10'd49: pixel <= 24'h75_B8_FF;
                10'd50: pixel <= 24'hB8_FF_50;
                10'd51: pixel <= 24'hFF_52_74;
                10'd52: pixel <= 24'h54_74_B6;
                10'd53: pixel <= 24'h75_B6_FF;
                10'd54: pixel <= 24'hB5_FF_52;
                10'd55: pixel <= 24'hFF_51_74;
                10'd56: pixel <= 24'h51_73_B7;
                10'd57: pixel <= 24'h74_B8_FF;
                10'd58: pixel <= 24'hB8_FF_52;
                10'd59: pixel <= 24'hFF_50_75;
                10'd60: pixel <= 24'h52_74_B8;
                10'd61: pixel <= 24'h73_B7_FF;
                10'd62: pixel <= 24'hB7_FF_51;
                10'd63: pixel <= 24'hFF_50_74;
                10'd64: pixel <= 24'h51_73_B7;
                10'd65: pixel <= 24'h74_B7_FF;
                10'd66: pixel <= 24'hB8_FF_4F;
                10'd67: pixel <= 24'hFF_52_74;
                10'd68: pixel <= 24'h50_75_B8;
                10'd69: pixel <= 24'h75_B8_FF;
                10'd70: pixel <= 24'hB7_FF_50;
                10'd71: pixel <= 24'hFF_4F_74;
                10'd72: pixel <= 24'h51_73_B9;
                10'd73: pixel <= 24'h74_B9_FF;
                10'd74: pixel <= 24'hB9_FF_4F;
                10'd75: pixel <= 24'hFF_51_73;
                10'd76: pixel <= 24'h51_73_B9;
                10'd77: pixel <= 24'h74_B5_FF;
                10'd78: pixel <= 24'hB4_FF_51;
                10'd79: pixel <= 24'hFF_52_75;
                10'd80: pixel <= 24'h50_76_B6;
                10'd81: pixel <= 24'h76_B8_FF;
                10'd82: pixel <= 24'hB8_FF_4F;
                10'd83: pixel <= 24'hFF_4F_76;
                10'd84: pixel <= 24'h50_75_B8;
                10'd85: pixel <= 24'h75_B8_FF;
                10'd86: pixel <= 24'hB6_FF_50;
                10'd87: pixel <= 24'hFF_50_76;
                10'd88: pixel <= 24'h52_7A_BC;
                10'd89: pixel <= 24'h7A_BC_FF;
                10'd90: pixel <= 24'hBA_FF_52;
                10'd91: pixel <= 24'hFF_54_79;
                10'd92: pixel <= 24'h40_55_AA;
                10'd93: pixel <= 24'h00_00_0C;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd65: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'hAA_00_00;
                10'd7: pixel <= 24'h0C_40_55;
                10'd8: pixel <= 24'h57_79_BD;
                10'd9: pixel <= 24'h7A_BC_FF;
                10'd10: pixel <= 24'hBC_FF_52;
                10'd11: pixel <= 24'hFF_52_7A;
                10'd12: pixel <= 24'h52_7A_BC;
                10'd13: pixel <= 24'h7A_BC_FF;
                10'd14: pixel <= 24'hBC_FF_52;
                10'd15: pixel <= 24'hFF_52_7A;
                10'd16: pixel <= 24'h52_7A_BC;
                10'd17: pixel <= 24'h7A_BC_FF;
                10'd18: pixel <= 24'hBC_FF_52;
                10'd19: pixel <= 24'hFF_52_7A;
                10'd20: pixel <= 24'h52_7A_BC;
                10'd21: pixel <= 24'h7A_BC_FF;
                10'd22: pixel <= 24'hBC_FF_52;
                10'd23: pixel <= 24'hFF_52_7A;
                10'd24: pixel <= 24'h52_7A_BC;
                10'd25: pixel <= 24'h7A_BC_FF;
                10'd26: pixel <= 24'hBC_FF_52;
                10'd27: pixel <= 24'hFF_52_7A;
                10'd28: pixel <= 24'h52_7A_BC;
                10'd29: pixel <= 24'h7A_BC_FF;
                10'd30: pixel <= 24'hBC_FF_52;
                10'd31: pixel <= 24'hFF_52_7A;
                10'd32: pixel <= 24'h52_7A_BC;
                10'd33: pixel <= 24'h7A_BC_FF;
                10'd34: pixel <= 24'hBC_FF_52;
                10'd35: pixel <= 24'hFF_52_7A;
                10'd36: pixel <= 24'h52_7A_BC;
                10'd37: pixel <= 24'h7A_BC_FF;
                10'd38: pixel <= 24'hBC_FF_52;
                10'd39: pixel <= 24'hFF_52_7A;
                10'd40: pixel <= 24'h52_7A_BC;
                10'd41: pixel <= 24'h7A_BC_FF;
                10'd42: pixel <= 24'hBC_FF_52;
                10'd43: pixel <= 24'hFF_52_7A;
                10'd44: pixel <= 24'h52_7A_BC;
                10'd45: pixel <= 24'h7A_BC_FF;
                10'd46: pixel <= 24'hBC_FF_52;
                10'd47: pixel <= 24'hFF_52_7A;
                10'd48: pixel <= 24'h52_7A_BC;
                10'd49: pixel <= 24'h7A_BC_FF;
                10'd50: pixel <= 24'hBC_FF_52;
                10'd51: pixel <= 24'hFF_52_7A;
                10'd52: pixel <= 24'h52_7A_BC;
                10'd53: pixel <= 24'h7A_BC_FF;
                10'd54: pixel <= 24'hBC_FF_52;
                10'd55: pixel <= 24'hFF_52_7A;
                10'd56: pixel <= 24'h52_7A_BC;
                10'd57: pixel <= 24'h79_BA_FF;
                10'd58: pixel <= 24'hAA_FF_54;
                10'd59: pixel <= 24'h0C_40_55;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd66: case (x)
                10'd0: pixel <= 24'h54_7B_BD;
                10'd1: pixel <= 24'h7A_BD_FF;
                10'd2: pixel <= 24'hBD_FF_55;
                10'd3: pixel <= 24'hFF_55_7A;
                10'd4: pixel <= 24'h55_7A_BD;
                10'd5: pixel <= 24'h7A_BD_FF;
                10'd6: pixel <= 24'hBD_FF_55;
                10'd7: pixel <= 24'hFF_55_7A;
                10'd8: pixel <= 24'h55_7A_BD;
                10'd9: pixel <= 24'h7B_BD_FF;
                10'd10: pixel <= 24'hBD_FF_54;
                10'd11: pixel <= 24'hFF_55_7A;
                10'd12: pixel <= 24'h54_7B_BD;
                10'd13: pixel <= 24'h7A_BD_FF;
                10'd14: pixel <= 24'hBD_FF_55;
                10'd15: pixel <= 24'hFF_55_7A;
                10'd16: pixel <= 24'h55_7A_BD;
                10'd17: pixel <= 24'h7A_BD_FF;
                10'd18: pixel <= 24'hBD_FF_55;
                10'd19: pixel <= 24'hFF_54_7B;
                10'd20: pixel <= 24'h55_7A_BD;
                10'd21: pixel <= 24'h7B_BD_FF;
                10'd22: pixel <= 24'hBD_FF_54;
                10'd23: pixel <= 24'hFF_55_7A;
                10'd24: pixel <= 24'h57_7A_BB;
                10'd25: pixel <= 24'h55_AA_FF;
                10'd26: pixel <= 24'h00_0C_40;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h00_00_00;
                10'd74: pixel <= 24'h00_00_00;
                10'd75: pixel <= 24'h00_00_00;
                10'd76: pixel <= 24'h00_00_00;
                10'd77: pixel <= 24'h00_00_00;
                10'd78: pixel <= 24'h00_00_00;
                10'd79: pixel <= 24'h00_00_00;
                10'd80: pixel <= 24'h00_00_00;
                10'd81: pixel <= 24'h00_00_00;
                10'd82: pixel <= 24'h00_00_00;
                10'd83: pixel <= 24'h00_00_00;
                10'd84: pixel <= 24'h00_00_00;
                10'd85: pixel <= 24'h00_00_00;
                10'd86: pixel <= 24'h00_00_00;
                10'd87: pixel <= 24'h00_00_00;
                10'd88: pixel <= 24'h00_00_00;
                10'd89: pixel <= 24'h00_00_00;
                10'd90: pixel <= 24'h00_00_00;
                10'd91: pixel <= 24'h00_00_00;
                10'd92: pixel <= 24'h00_00_00;
                10'd93: pixel <= 24'h00_00_00;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
            10'd67: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h00_00_00;
                10'd41: pixel <= 24'h00_00_00;
                10'd42: pixel <= 24'h00_00_00;
                10'd43: pixel <= 24'h00_00_00;
                10'd44: pixel <= 24'h00_00_00;
                10'd45: pixel <= 24'h00_00_00;
                10'd46: pixel <= 24'h00_00_00;
                10'd47: pixel <= 24'h00_00_00;
                10'd48: pixel <= 24'h00_00_00;
                10'd49: pixel <= 24'h00_00_00;
                10'd50: pixel <= 24'h00_00_00;
                10'd51: pixel <= 24'h00_00_00;
                10'd52: pixel <= 24'h00_00_00;
                10'd53: pixel <= 24'h00_00_00;
                10'd54: pixel <= 24'h00_00_00;
                10'd55: pixel <= 24'h00_00_00;
                10'd56: pixel <= 24'h00_00_00;
                10'd57: pixel <= 24'h00_00_00;
                10'd58: pixel <= 24'h00_00_00;
                10'd59: pixel <= 24'h00_00_00;
                10'd60: pixel <= 24'h00_00_00;
                10'd61: pixel <= 24'h00_00_00;
                10'd62: pixel <= 24'h00_00_00;
                10'd63: pixel <= 24'h00_00_00;
                10'd64: pixel <= 24'h00_00_00;
                10'd65: pixel <= 24'h00_00_00;
                10'd66: pixel <= 24'h00_00_00;
                10'd67: pixel <= 24'h00_00_00;
                10'd68: pixel <= 24'h00_00_00;
                10'd69: pixel <= 24'h00_00_00;
                10'd70: pixel <= 24'h00_00_00;
                10'd71: pixel <= 24'h00_00_00;
                10'd72: pixel <= 24'h00_00_00;
                10'd73: pixel <= 24'h55_AA_00;
                10'd74: pixel <= 24'hBD_0C_40;
                10'd75: pixel <= 24'hFF_57_79;
                10'd76: pixel <= 24'h54_7B_BD;
                10'd77: pixel <= 24'h7A_BD_FF;
                10'd78: pixel <= 24'hBD_FF_55;
                10'd79: pixel <= 24'hFF_54_7B;
                10'd80: pixel <= 24'h55_7A_BD;
                10'd81: pixel <= 24'h7A_BD_FF;
                10'd82: pixel <= 24'hBD_FF_55;
                10'd83: pixel <= 24'hFF_54_7B;
                10'd84: pixel <= 24'h55_7A_BD;
                10'd85: pixel <= 24'h7A_BD_FF;
                10'd86: pixel <= 24'hBD_FF_55;
                10'd87: pixel <= 24'hFF_55_7A;
                10'd88: pixel <= 24'h54_7B_BD;
                10'd89: pixel <= 24'h7A_BD_FF;
                10'd90: pixel <= 24'hBD_FF_55;
                10'd91: pixel <= 24'hFF_54_7B;
                10'd92: pixel <= 24'h55_7A_BD;
                10'd93: pixel <= 24'h7A_BD_FF;
                10'd94: pixel <= 24'hBD_FF_55;
                10'd95: pixel <= 24'hFF_55_7A;
                10'd96: pixel <= 24'h55_7A_BD;
                10'd97: pixel <= 24'h7B_BD_FF;
                10'd98: pixel <= 24'hBD_FF_54;
                10'd99: pixel <= 24'hFF_55_7A;
            endcase
            10'd68: case (x)
                10'd0: pixel <= 24'h00_00_00;
                10'd1: pixel <= 24'h00_00_00;
                10'd2: pixel <= 24'h00_00_00;
                10'd3: pixel <= 24'h00_00_00;
                10'd4: pixel <= 24'h00_00_00;
                10'd5: pixel <= 24'h00_00_00;
                10'd6: pixel <= 24'h00_00_00;
                10'd7: pixel <= 24'h00_00_00;
                10'd8: pixel <= 24'h00_00_00;
                10'd9: pixel <= 24'h00_00_00;
                10'd10: pixel <= 24'h00_00_00;
                10'd11: pixel <= 24'h00_00_00;
                10'd12: pixel <= 24'h00_00_00;
                10'd13: pixel <= 24'h00_00_00;
                10'd14: pixel <= 24'h00_00_00;
                10'd15: pixel <= 24'h00_00_00;
                10'd16: pixel <= 24'h00_00_00;
                10'd17: pixel <= 24'h00_00_00;
                10'd18: pixel <= 24'h00_00_00;
                10'd19: pixel <= 24'h00_00_00;
                10'd20: pixel <= 24'h00_00_00;
                10'd21: pixel <= 24'h00_00_00;
                10'd22: pixel <= 24'h00_00_00;
                10'd23: pixel <= 24'h00_00_00;
                10'd24: pixel <= 24'h00_00_00;
                10'd25: pixel <= 24'h00_00_00;
                10'd26: pixel <= 24'h00_00_00;
                10'd27: pixel <= 24'h00_00_00;
                10'd28: pixel <= 24'h00_00_00;
                10'd29: pixel <= 24'h00_00_00;
                10'd30: pixel <= 24'h00_00_00;
                10'd31: pixel <= 24'h00_00_00;
                10'd32: pixel <= 24'h00_00_00;
                10'd33: pixel <= 24'h00_00_00;
                10'd34: pixel <= 24'h00_00_00;
                10'd35: pixel <= 24'h00_00_00;
                10'd36: pixel <= 24'h00_00_00;
                10'd37: pixel <= 24'h00_00_00;
                10'd38: pixel <= 24'h00_00_00;
                10'd39: pixel <= 24'h00_00_00;
                10'd40: pixel <= 24'h40_55_AA;
                10'd41: pixel <= 24'h42_83_0C;
                10'd42: pixel <= 24'h85_FF_1F;
                10'd43: pixel <= 24'hFF_22_42;
                10'd44: pixel <= 24'h22_42_85;
                10'd45: pixel <= 24'h41_85_FF;
                10'd46: pixel <= 24'h85_FF_23;
                10'd47: pixel <= 24'hFF_22_42;
                10'd48: pixel <= 24'h22_42_85;
                10'd49: pixel <= 24'h43_85_FF;
                10'd50: pixel <= 24'h85_FF_20;
                10'd51: pixel <= 24'hFF_22_42;
                10'd52: pixel <= 24'h22_42_85;
                10'd53: pixel <= 24'h42_85_FF;
                10'd54: pixel <= 24'h85_FF_22;
                10'd55: pixel <= 24'hFF_23_41;
                10'd56: pixel <= 24'h22_42_85;
                10'd57: pixel <= 24'h42_85_FF;
                10'd58: pixel <= 24'h85_FF_22;
                10'd59: pixel <= 24'hFF_22_42;
                10'd60: pixel <= 24'h22_42_85;
                10'd61: pixel <= 24'h42_85_FF;
                10'd62: pixel <= 24'h85_FF_22;
                10'd63: pixel <= 24'hFF_22_42;
                10'd64: pixel <= 24'h22_42_85;
                10'd65: pixel <= 24'h42_85_FF;
                10'd66: pixel <= 24'h85_FF_22;
                10'd67: pixel <= 24'hFF_23_41;
                10'd68: pixel <= 24'h22_42_85;
                10'd69: pixel <= 24'h42_85_FF;
                10'd70: pixel <= 24'h85_FF_22;
                10'd71: pixel <= 24'hFF_22_42;
                10'd72: pixel <= 24'h22_42_85;
                10'd73: pixel <= 24'h42_85_FF;
                10'd74: pixel <= 24'h85_FF_22;
                10'd75: pixel <= 24'hFF_22_42;
                10'd76: pixel <= 24'h23_41_85;
                10'd77: pixel <= 24'h42_85_FF;
                10'd78: pixel <= 24'h85_FF_22;
                10'd79: pixel <= 24'hFF_22_42;
                10'd80: pixel <= 24'h22_42_85;
                10'd81: pixel <= 24'h42_85_FF;
                10'd82: pixel <= 24'h85_FF_22;
                10'd83: pixel <= 24'hFF_22_42;
                10'd84: pixel <= 24'h22_42_85;
                10'd85: pixel <= 24'h42_85_FF;
                10'd86: pixel <= 24'h85_FF_22;
                10'd87: pixel <= 24'hFF_22_42;
                10'd88: pixel <= 24'h23_41_85;
                10'd89: pixel <= 24'h42_85_FF;
                10'd90: pixel <= 24'h83_FF_22;
                10'd91: pixel <= 24'hFF_22_43;
                10'd92: pixel <= 24'h40_55_AA;
                10'd93: pixel <= 24'h00_00_0C;
                10'd94: pixel <= 24'h00_00_00;
                10'd95: pixel <= 24'h00_00_00;
                10'd96: pixel <= 24'h00_00_00;
                10'd97: pixel <= 24'h00_00_00;
                10'd98: pixel <= 24'h00_00_00;
                10'd99: pixel <= 24'h00_00_00;
            endcase
        endcase

        end

endmodule
